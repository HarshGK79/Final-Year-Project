VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ALU
  CLASS BLOCK ;
  FOREIGN ALU ;
  ORIGIN 2.600 3.000 ;
  SIZE 103.600 BY 86.200 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.200 80.200 98.200 80.800 ;
        RECT 1.400 76.500 1.800 80.200 ;
        RECT 3.800 77.900 4.200 80.200 ;
        RECT 4.600 77.900 5.000 80.200 ;
        RECT 6.200 77.900 6.600 80.200 ;
        RECT 7.800 77.900 8.200 80.200 ;
        RECT 8.600 77.900 9.000 80.200 ;
        RECT 10.200 77.900 10.600 80.200 ;
        RECT 11.000 77.900 11.400 80.200 ;
        RECT 14.200 75.900 14.600 80.200 ;
        RECT 15.000 77.900 15.400 80.200 ;
        RECT 16.600 77.900 17.000 80.200 ;
        RECT 17.400 75.900 17.800 80.200 ;
        RECT 19.800 77.900 20.200 80.200 ;
        RECT 21.400 77.900 21.800 80.200 ;
        RECT 23.000 76.100 23.400 80.200 ;
        RECT 24.600 77.900 25.000 80.200 ;
        RECT 25.400 77.900 25.800 80.200 ;
        RECT 27.000 77.900 27.400 80.200 ;
        RECT 30.200 77.900 30.600 80.200 ;
        RECT 31.800 75.900 32.200 80.200 ;
        RECT 34.200 75.900 34.600 80.200 ;
        RECT 35.800 75.900 36.200 80.200 ;
        RECT 36.600 77.900 37.000 80.200 ;
        RECT 38.200 78.100 38.600 80.200 ;
        RECT 41.400 76.500 41.800 80.200 ;
        RECT 43.800 77.900 44.200 80.200 ;
        RECT 44.600 75.900 45.000 80.200 ;
        RECT 47.800 75.900 48.200 80.200 ;
        RECT 48.600 75.900 49.000 80.200 ;
        RECT 52.600 75.900 53.000 80.200 ;
        RECT 53.400 75.900 53.800 80.200 ;
        RECT 55.000 75.900 55.400 80.200 ;
        RECT 60.600 76.900 61.000 80.200 ;
        RECT 63.800 76.500 64.200 80.200 ;
        RECT 65.700 77.900 66.100 80.200 ;
        RECT 67.800 75.900 68.200 80.200 ;
        RECT 70.200 77.900 70.600 80.200 ;
        RECT 71.800 78.100 72.200 80.200 ;
        RECT 74.200 77.900 74.600 80.200 ;
        RECT 75.800 78.100 76.200 80.200 ;
        RECT 77.400 77.900 77.800 80.200 ;
        RECT 79.000 76.500 79.400 80.200 ;
        RECT 82.200 76.900 82.600 80.200 ;
        RECT 88.600 76.500 89.000 80.200 ;
        RECT 91.000 76.500 91.400 80.200 ;
        RECT 93.400 76.500 93.800 80.200 ;
        RECT 95.800 76.500 96.200 80.200 ;
        RECT 5.400 60.800 5.800 64.100 ;
        RECT 7.000 60.800 7.400 63.100 ;
        RECT 8.600 60.800 9.000 63.100 ;
        RECT 11.000 60.800 11.400 65.100 ;
        RECT 12.600 60.800 13.000 62.900 ;
        RECT 14.200 60.800 14.600 63.100 ;
        RECT 15.000 60.800 15.400 63.100 ;
        RECT 16.600 60.800 17.000 63.100 ;
        RECT 17.400 60.800 17.800 63.100 ;
        RECT 19.000 60.800 19.400 63.100 ;
        RECT 19.800 60.800 20.200 65.100 ;
        RECT 23.800 60.800 24.200 65.100 ;
        RECT 24.600 60.800 25.000 65.100 ;
        RECT 28.600 60.800 29.000 65.100 ;
        RECT 31.000 60.800 31.400 65.100 ;
        RECT 33.400 60.800 33.800 65.100 ;
        RECT 35.800 60.800 36.200 65.100 ;
        RECT 39.800 60.800 40.200 65.100 ;
        RECT 40.600 60.800 41.000 65.100 ;
        RECT 43.000 60.800 43.400 65.100 ;
        RECT 47.000 60.800 47.400 64.500 ;
        RECT 48.900 60.800 49.300 63.100 ;
        RECT 51.000 60.800 51.400 65.100 ;
        RECT 51.800 60.800 52.200 65.100 ;
        RECT 55.000 60.800 55.400 64.500 ;
        RECT 56.900 60.800 57.300 63.100 ;
        RECT 59.000 60.800 59.400 65.100 ;
        RECT 59.800 60.800 60.200 65.100 ;
        RECT 63.000 60.800 63.400 65.100 ;
        RECT 63.800 60.800 64.200 65.100 ;
        RECT 66.200 60.800 66.600 65.100 ;
        RECT 69.400 60.800 69.800 63.100 ;
        RECT 71.000 60.800 71.400 62.900 ;
        RECT 72.600 60.800 73.000 63.100 ;
        RECT 74.200 60.800 74.600 63.100 ;
        RECT 75.000 60.800 75.400 65.100 ;
        RECT 77.100 60.800 77.500 63.100 ;
        RECT 78.200 60.800 78.600 65.100 ;
        RECT 80.600 60.800 81.000 65.100 ;
        RECT 83.800 60.800 84.200 62.900 ;
        RECT 85.400 60.800 85.800 63.100 ;
        RECT 87.800 60.800 88.200 64.500 ;
        RECT 91.000 60.800 91.400 64.500 ;
        RECT 93.400 60.800 93.800 63.100 ;
        RECT 94.200 60.800 94.600 63.100 ;
        RECT 95.800 60.800 96.200 63.100 ;
        RECT 0.200 60.200 98.200 60.800 ;
        RECT 0.600 57.900 1.000 60.200 ;
        RECT 2.200 57.900 2.600 60.200 ;
        RECT 3.000 57.900 3.400 60.200 ;
        RECT 4.600 58.100 5.000 60.200 ;
        RECT 6.200 57.900 6.600 60.200 ;
        RECT 7.800 56.100 8.200 60.200 ;
        RECT 9.400 55.900 9.800 60.200 ;
        RECT 12.600 55.900 13.000 60.200 ;
        RECT 13.400 57.900 13.800 60.200 ;
        RECT 15.000 57.900 15.400 60.200 ;
        RECT 15.800 55.900 16.200 60.200 ;
        RECT 17.400 55.900 17.800 60.200 ;
        RECT 19.500 57.900 19.900 60.200 ;
        RECT 20.600 57.900 21.000 60.200 ;
        RECT 22.200 58.100 22.600 60.200 ;
        RECT 24.100 57.900 24.500 60.200 ;
        RECT 26.200 55.900 26.600 60.200 ;
        RECT 30.200 55.900 30.600 60.200 ;
        RECT 31.000 57.900 31.400 60.200 ;
        RECT 32.600 57.900 33.000 60.200 ;
        RECT 33.400 57.900 33.800 60.200 ;
        RECT 35.800 56.500 36.200 60.200 ;
        RECT 39.300 57.900 39.700 60.200 ;
        RECT 41.400 55.900 41.800 60.200 ;
        RECT 43.800 55.900 44.200 60.200 ;
        RECT 44.900 57.900 45.300 60.200 ;
        RECT 47.000 55.900 47.400 60.200 ;
        RECT 47.800 57.900 48.200 60.200 ;
        RECT 49.400 57.900 49.800 60.200 ;
        RECT 51.000 57.900 51.400 60.200 ;
        RECT 52.100 57.900 52.500 60.200 ;
        RECT 54.200 55.900 54.600 60.200 ;
        RECT 55.300 57.900 55.700 60.200 ;
        RECT 57.400 55.900 57.800 60.200 ;
        RECT 59.800 55.900 60.200 60.200 ;
        RECT 60.600 55.900 61.000 60.200 ;
        RECT 63.800 55.900 64.200 60.200 ;
        RECT 65.400 57.900 65.800 60.200 ;
        RECT 66.200 55.900 66.600 60.200 ;
        RECT 71.800 55.900 72.200 60.200 ;
        RECT 72.600 57.900 73.000 60.200 ;
        RECT 74.200 58.100 74.600 60.200 ;
        RECT 75.800 55.900 76.200 60.200 ;
        RECT 78.200 55.900 78.600 60.200 ;
        RECT 80.900 57.900 81.300 60.200 ;
        RECT 83.000 55.900 83.400 60.200 ;
        RECT 85.400 55.900 85.800 60.200 ;
        RECT 86.500 57.900 86.900 60.200 ;
        RECT 88.600 55.900 89.000 60.200 ;
        RECT 90.200 57.900 90.600 60.200 ;
        RECT 91.800 55.900 92.200 60.200 ;
        RECT 93.400 56.500 93.800 60.200 ;
        RECT 95.000 55.900 95.400 60.200 ;
        RECT 97.100 57.900 97.500 60.200 ;
        RECT 0.600 40.800 1.000 45.100 ;
        RECT 2.200 40.800 2.600 43.100 ;
        RECT 3.800 40.800 4.200 43.100 ;
        RECT 4.600 40.800 5.000 45.100 ;
        RECT 6.700 40.800 7.100 43.100 ;
        RECT 7.800 40.800 8.200 43.100 ;
        RECT 9.400 40.800 9.800 44.900 ;
        RECT 12.600 40.800 13.000 45.100 ;
        RECT 15.000 40.800 15.400 44.500 ;
        RECT 17.700 40.800 18.100 45.100 ;
        RECT 19.800 40.800 20.200 45.100 ;
        RECT 21.900 40.800 22.300 43.100 ;
        RECT 23.000 40.800 23.400 43.100 ;
        RECT 24.600 40.800 25.000 42.900 ;
        RECT 26.200 40.800 26.600 43.100 ;
        RECT 27.800 40.800 28.200 43.100 ;
        RECT 30.200 40.800 30.600 43.100 ;
        RECT 31.800 40.800 32.200 43.100 ;
        RECT 35.000 40.800 35.400 44.500 ;
        RECT 36.600 40.800 37.000 43.100 ;
        RECT 38.200 40.800 38.600 43.100 ;
        RECT 41.400 40.800 41.800 44.500 ;
        RECT 43.300 40.800 43.700 43.100 ;
        RECT 45.400 40.800 45.800 45.100 ;
        RECT 46.200 40.800 46.600 45.100 ;
        RECT 48.600 40.800 49.000 45.100 ;
        RECT 51.000 40.800 51.400 45.100 ;
        RECT 52.100 40.800 52.500 43.100 ;
        RECT 54.200 40.800 54.600 45.100 ;
        RECT 56.600 40.800 57.000 44.500 ;
        RECT 58.200 40.800 58.600 43.100 ;
        RECT 59.800 40.800 60.200 42.900 ;
        RECT 61.400 40.800 61.800 45.100 ;
        RECT 63.500 40.800 63.900 43.100 ;
        RECT 64.600 40.800 65.000 45.100 ;
        RECT 66.700 40.800 67.100 43.100 ;
        RECT 70.200 40.800 70.600 44.500 ;
        RECT 72.600 40.800 73.000 43.100 ;
        RECT 74.200 40.800 74.600 42.900 ;
        RECT 75.800 40.800 76.200 45.100 ;
        RECT 77.400 40.800 77.800 45.100 ;
        RECT 79.500 40.800 79.900 43.100 ;
        RECT 81.400 40.800 81.800 44.500 ;
        RECT 83.800 40.800 84.200 45.100 ;
        RECT 91.000 40.800 91.400 44.100 ;
        RECT 93.400 40.800 93.800 44.500 ;
        RECT 95.000 40.800 95.400 43.100 ;
        RECT 96.600 40.800 97.000 44.900 ;
        RECT 0.200 40.200 98.200 40.800 ;
        RECT 0.600 35.900 1.000 40.200 ;
        RECT 2.700 37.900 3.100 40.200 ;
        RECT 4.600 36.500 5.000 40.200 ;
        RECT 7.800 35.900 8.200 40.200 ;
        RECT 9.400 35.900 9.800 40.200 ;
        RECT 11.500 37.900 11.900 40.200 ;
        RECT 12.600 35.900 13.000 40.200 ;
        RECT 16.300 35.900 16.700 40.200 ;
        RECT 19.000 36.500 19.400 40.200 ;
        RECT 22.200 36.500 22.600 40.200 ;
        RECT 26.200 35.900 26.600 40.200 ;
        RECT 28.600 35.900 29.000 40.200 ;
        RECT 30.700 37.900 31.100 40.200 ;
        RECT 31.800 37.900 32.200 40.200 ;
        RECT 33.400 37.900 33.800 40.200 ;
        RECT 35.000 36.500 35.400 40.200 ;
        RECT 37.400 35.900 37.800 40.200 ;
        RECT 39.500 37.900 39.900 40.200 ;
        RECT 41.400 37.900 41.800 40.200 ;
        RECT 42.200 35.900 42.600 40.200 ;
        RECT 44.600 35.900 45.000 40.200 ;
        RECT 46.700 37.900 47.100 40.200 ;
        RECT 49.400 35.900 49.800 40.200 ;
        RECT 51.000 36.500 51.400 40.200 ;
        RECT 54.500 37.900 54.900 40.200 ;
        RECT 56.600 35.900 57.000 40.200 ;
        RECT 58.200 37.900 58.600 40.200 ;
        RECT 63.800 36.900 64.200 40.200 ;
        RECT 65.400 35.900 65.800 40.200 ;
        RECT 67.500 37.900 67.900 40.200 ;
        RECT 70.500 37.900 70.900 40.200 ;
        RECT 72.600 35.900 73.000 40.200 ;
        RECT 73.400 37.900 73.800 40.200 ;
        RECT 75.000 37.900 75.400 40.200 ;
        RECT 75.800 35.900 76.200 40.200 ;
        RECT 77.900 37.900 78.300 40.200 ;
        RECT 79.000 37.900 79.400 40.200 ;
        RECT 80.900 37.900 81.300 40.200 ;
        RECT 83.000 35.900 83.400 40.200 ;
        RECT 84.100 37.900 84.500 40.200 ;
        RECT 86.200 35.900 86.600 40.200 ;
        RECT 87.800 35.900 88.200 40.200 ;
        RECT 88.600 35.900 89.000 40.200 ;
        RECT 90.700 37.900 91.100 40.200 ;
        RECT 91.800 37.900 92.200 40.200 ;
        RECT 93.400 37.900 93.800 40.200 ;
        RECT 95.000 37.900 95.400 40.200 ;
        RECT 1.400 20.800 1.800 24.500 ;
        RECT 3.000 20.800 3.400 23.100 ;
        RECT 4.600 20.800 5.000 23.100 ;
        RECT 6.200 20.800 6.600 22.900 ;
        RECT 7.800 20.800 8.200 23.100 ;
        RECT 8.900 20.800 9.300 23.100 ;
        RECT 11.000 20.800 11.400 25.100 ;
        RECT 16.600 20.800 17.000 24.100 ;
        RECT 18.500 20.800 18.900 23.100 ;
        RECT 20.600 20.800 21.000 25.100 ;
        RECT 21.700 20.800 22.100 23.100 ;
        RECT 23.800 20.800 24.200 25.100 ;
        RECT 25.900 20.800 26.300 25.100 ;
        RECT 31.000 20.800 31.400 25.100 ;
        RECT 31.800 20.800 32.200 23.100 ;
        RECT 33.400 20.800 33.800 22.900 ;
        RECT 35.000 20.800 35.400 25.100 ;
        RECT 37.100 20.800 37.500 23.100 ;
        RECT 39.000 20.800 39.400 23.100 ;
        RECT 39.800 20.800 40.200 25.100 ;
        RECT 42.200 20.800 42.600 25.100 ;
        RECT 44.300 20.800 44.700 23.100 ;
        RECT 46.200 20.800 46.600 23.100 ;
        RECT 47.800 20.800 48.200 24.500 ;
        RECT 51.000 20.800 51.400 23.100 ;
        RECT 55.000 20.800 55.400 24.500 ;
        RECT 57.400 20.800 57.800 24.500 ;
        RECT 60.600 20.800 61.000 24.500 ;
        RECT 63.000 20.800 63.400 25.100 ;
        RECT 65.100 20.800 65.500 23.100 ;
        RECT 67.800 20.800 68.200 25.100 ;
        RECT 70.500 20.800 70.900 23.100 ;
        RECT 72.600 20.800 73.000 25.100 ;
        RECT 73.400 20.800 73.800 23.100 ;
        RECT 75.000 20.800 75.400 23.100 ;
        RECT 76.100 20.800 76.500 23.100 ;
        RECT 78.200 20.800 78.600 25.100 ;
        RECT 80.600 20.800 81.000 25.100 ;
        RECT 82.200 20.800 82.600 24.500 ;
        RECT 84.900 20.800 85.300 23.100 ;
        RECT 87.000 20.800 87.400 25.100 ;
        RECT 88.600 20.800 89.000 25.100 ;
        RECT 89.400 20.800 89.800 23.100 ;
        RECT 91.000 20.800 91.400 23.100 ;
        RECT 93.400 20.800 93.800 25.100 ;
        RECT 94.500 20.800 94.900 23.100 ;
        RECT 96.600 20.800 97.000 25.100 ;
        RECT 0.200 20.200 98.200 20.800 ;
        RECT 5.400 16.900 5.800 20.200 ;
        RECT 7.000 15.900 7.400 20.200 ;
        RECT 9.100 17.900 9.500 20.200 ;
        RECT 11.000 18.100 11.400 20.200 ;
        RECT 12.600 17.900 13.000 20.200 ;
        RECT 13.400 17.900 13.800 20.200 ;
        RECT 15.000 17.900 15.400 20.200 ;
        RECT 15.800 17.900 16.200 20.200 ;
        RECT 17.400 17.900 17.800 20.200 ;
        RECT 19.000 16.500 19.400 20.200 ;
        RECT 21.700 17.900 22.100 20.200 ;
        RECT 23.800 15.900 24.200 20.200 ;
        RECT 24.600 17.900 25.000 20.200 ;
        RECT 26.200 17.900 26.600 20.200 ;
        RECT 28.600 17.900 29.000 20.200 ;
        RECT 30.200 17.900 30.600 20.200 ;
        RECT 31.000 17.900 31.400 20.200 ;
        RECT 32.600 18.100 33.000 20.200 ;
        RECT 34.200 15.900 34.600 20.200 ;
        RECT 36.300 17.900 36.700 20.200 ;
        RECT 37.400 15.900 37.800 20.200 ;
        RECT 41.400 16.500 41.800 20.200 ;
        RECT 43.800 16.500 44.200 20.200 ;
        RECT 47.000 18.100 47.400 20.200 ;
        RECT 48.600 17.900 49.000 20.200 ;
        RECT 51.800 16.500 52.200 20.200 ;
        RECT 53.400 15.900 53.800 20.200 ;
        RECT 55.500 17.900 55.900 20.200 ;
        RECT 57.400 16.900 57.800 20.200 ;
        RECT 63.000 15.900 63.400 20.200 ;
        RECT 65.100 17.900 65.500 20.200 ;
        RECT 66.500 17.900 66.900 20.200 ;
        RECT 68.600 15.900 69.000 20.200 ;
        RECT 71.000 15.900 71.400 20.200 ;
        RECT 72.600 15.900 73.000 20.200 ;
        RECT 75.800 15.900 76.200 20.200 ;
        RECT 77.400 16.500 77.800 20.200 ;
        RECT 80.100 17.900 80.500 20.200 ;
        RECT 82.200 15.900 82.600 20.200 ;
        RECT 83.000 15.900 83.400 20.200 ;
        RECT 85.100 17.900 85.500 20.200 ;
        RECT 87.800 16.500 88.200 20.200 ;
        RECT 89.400 17.900 89.800 20.200 ;
        RECT 91.000 18.100 91.400 20.200 ;
        RECT 94.200 16.500 94.600 20.200 ;
        RECT 1.400 0.800 1.900 4.400 ;
        RECT 4.500 1.100 5.000 4.400 ;
        RECT 4.500 0.800 4.900 1.100 ;
        RECT 6.200 0.800 6.600 3.100 ;
        RECT 7.800 0.800 8.200 4.900 ;
        RECT 10.700 0.800 11.100 5.100 ;
        RECT 12.600 0.800 13.000 3.100 ;
        RECT 14.200 0.800 14.600 3.100 ;
        RECT 15.800 0.800 16.200 4.500 ;
        RECT 19.000 0.800 19.400 3.100 ;
        RECT 20.600 0.800 21.000 3.100 ;
        RECT 23.000 0.800 23.400 5.100 ;
        RECT 23.800 0.800 24.200 5.100 ;
        RECT 27.000 0.800 27.400 5.100 ;
        RECT 31.000 0.800 31.400 5.100 ;
        RECT 31.800 0.800 32.200 5.100 ;
        RECT 33.900 0.800 34.300 3.100 ;
        RECT 35.000 0.800 35.400 3.100 ;
        RECT 36.600 0.800 37.000 3.100 ;
        RECT 38.500 0.800 38.900 5.100 ;
        RECT 41.400 0.800 41.800 4.500 ;
        RECT 45.400 0.800 45.800 4.900 ;
        RECT 47.000 0.800 47.400 3.100 ;
        RECT 48.600 1.100 49.100 4.400 ;
        RECT 48.700 0.800 49.100 1.100 ;
        RECT 51.700 0.800 52.200 4.400 ;
        RECT 54.200 0.800 54.600 4.500 ;
        RECT 56.600 0.800 57.000 4.500 ;
        RECT 59.000 0.800 59.500 4.400 ;
        RECT 62.100 1.100 62.600 4.400 ;
        RECT 62.100 0.800 62.500 1.100 ;
        RECT 66.200 0.800 66.600 4.500 ;
        RECT 69.400 0.800 69.800 3.100 ;
        RECT 71.000 0.800 71.400 3.100 ;
        RECT 71.800 0.800 72.200 5.100 ;
        RECT 73.400 0.800 73.800 3.100 ;
        RECT 75.000 0.800 75.400 3.100 ;
        RECT 75.800 0.800 76.200 3.100 ;
        RECT 77.400 0.800 77.800 5.100 ;
        RECT 79.500 0.800 79.900 3.100 ;
        RECT 81.400 0.800 81.800 5.100 ;
        RECT 82.200 0.800 82.600 3.100 ;
        RECT 83.800 0.800 84.200 3.100 ;
        RECT 86.200 0.800 86.600 5.100 ;
        RECT 87.800 0.800 88.200 4.500 ;
        RECT 90.200 0.800 90.600 3.100 ;
        RECT 91.800 0.800 92.300 4.400 ;
        RECT 94.900 1.100 95.400 4.400 ;
        RECT 94.900 0.800 95.300 1.100 ;
        RECT 0.200 0.200 98.200 0.800 ;
      LAYER via1 ;
        RECT 27.400 80.300 27.800 80.700 ;
        RECT 28.100 80.300 28.500 80.700 ;
        RECT 27.400 60.300 27.800 60.700 ;
        RECT 28.100 60.300 28.500 60.700 ;
        RECT 27.400 40.300 27.800 40.700 ;
        RECT 28.100 40.300 28.500 40.700 ;
        RECT 27.400 20.300 27.800 20.700 ;
        RECT 28.100 20.300 28.500 20.700 ;
        RECT 27.400 0.300 27.800 0.700 ;
        RECT 28.100 0.300 28.500 0.700 ;
      LAYER metal2 ;
        RECT 27.200 80.300 28.800 80.700 ;
        RECT 27.200 60.300 28.800 60.700 ;
        RECT 27.200 40.300 28.800 40.700 ;
        RECT 27.200 20.300 28.800 20.700 ;
        RECT 27.200 0.300 28.800 0.700 ;
      LAYER via2 ;
        RECT 27.400 80.300 27.800 80.700 ;
        RECT 28.100 80.300 28.500 80.700 ;
        RECT 27.400 60.300 27.800 60.700 ;
        RECT 28.100 60.300 28.500 60.700 ;
        RECT 27.400 40.300 27.800 40.700 ;
        RECT 28.100 40.300 28.500 40.700 ;
        RECT 27.400 20.300 27.800 20.700 ;
        RECT 28.100 20.300 28.500 20.700 ;
        RECT 27.400 0.300 27.800 0.700 ;
        RECT 28.100 0.300 28.500 0.700 ;
      LAYER metal3 ;
        RECT 27.200 80.300 28.800 80.700 ;
        RECT 27.200 60.300 28.800 60.700 ;
        RECT 27.200 40.300 28.800 40.700 ;
        RECT 27.200 20.300 28.800 20.700 ;
        RECT 27.200 0.300 28.800 0.700 ;
      LAYER via3 ;
        RECT 27.400 80.300 27.800 80.700 ;
        RECT 28.200 80.300 28.600 80.700 ;
        RECT 27.400 60.300 27.800 60.700 ;
        RECT 28.200 60.300 28.600 60.700 ;
        RECT 27.400 40.300 27.800 40.700 ;
        RECT 28.200 40.300 28.600 40.700 ;
        RECT 27.400 20.300 27.800 20.700 ;
        RECT 28.200 20.300 28.600 20.700 ;
        RECT 27.400 0.300 27.800 0.700 ;
        RECT 28.200 0.300 28.600 0.700 ;
      LAYER metal4 ;
        RECT 27.200 80.300 28.800 80.700 ;
        RECT 27.200 60.300 28.800 60.700 ;
        RECT 27.200 40.300 28.800 40.700 ;
        RECT 27.200 20.300 28.800 20.700 ;
        RECT 27.200 0.300 28.800 0.700 ;
      LAYER via4 ;
        RECT 27.400 80.300 27.800 80.700 ;
        RECT 28.100 80.300 28.500 80.700 ;
        RECT 27.400 60.300 27.800 60.700 ;
        RECT 28.100 60.300 28.500 60.700 ;
        RECT 27.400 40.300 27.800 40.700 ;
        RECT 28.100 40.300 28.500 40.700 ;
        RECT 27.400 20.300 27.800 20.700 ;
        RECT 28.100 20.300 28.500 20.700 ;
        RECT 27.400 0.300 27.800 0.700 ;
        RECT 28.100 0.300 28.500 0.700 ;
      LAYER metal5 ;
        RECT 27.200 80.200 28.800 80.700 ;
        RECT 27.200 60.200 28.800 60.700 ;
        RECT 27.200 40.200 28.800 40.700 ;
        RECT 27.200 20.200 28.800 20.700 ;
        RECT 27.200 0.200 28.800 0.700 ;
      LAYER via5 ;
        RECT 28.200 80.200 28.700 80.700 ;
        RECT 28.200 60.200 28.700 60.700 ;
        RECT 28.200 40.200 28.700 40.700 ;
        RECT 28.200 20.200 28.700 20.700 ;
        RECT 28.200 0.200 28.700 0.700 ;
      LAYER metal6 ;
        RECT 27.200 -3.000 28.800 83.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 1.400 70.800 1.800 73.100 ;
        RECT 3.800 70.800 4.200 72.100 ;
        RECT 4.600 70.800 5.000 72.100 ;
        RECT 7.800 70.800 8.200 73.100 ;
        RECT 8.600 70.800 9.000 73.100 ;
        RECT 11.000 70.800 11.400 72.100 ;
        RECT 12.600 70.800 13.000 72.100 ;
        RECT 14.200 70.800 14.600 72.100 ;
        RECT 15.000 70.800 15.400 73.100 ;
        RECT 17.400 70.800 17.800 72.100 ;
        RECT 19.000 70.800 19.400 72.100 ;
        RECT 19.800 70.800 20.200 73.100 ;
        RECT 23.300 70.800 23.700 73.000 ;
        RECT 25.400 70.800 25.800 73.100 ;
        RECT 30.200 70.800 30.600 72.100 ;
        RECT 31.800 70.800 32.200 73.100 ;
        RECT 32.600 70.800 33.000 72.100 ;
        RECT 34.200 70.800 34.600 72.100 ;
        RECT 35.800 70.800 36.200 73.100 ;
        RECT 36.600 70.800 37.000 74.100 ;
        RECT 39.800 70.800 40.200 72.100 ;
        RECT 41.900 70.800 42.300 73.100 ;
        RECT 43.800 70.800 44.200 72.100 ;
        RECT 44.600 70.800 45.000 72.100 ;
        RECT 46.200 70.800 46.600 72.100 ;
        RECT 47.800 70.800 48.200 73.100 ;
        RECT 48.600 70.800 49.000 72.100 ;
        RECT 50.200 70.800 50.600 72.100 ;
        RECT 51.000 70.800 51.400 72.100 ;
        RECT 52.600 70.800 53.000 72.100 ;
        RECT 53.400 70.800 53.800 73.100 ;
        RECT 55.000 70.800 55.400 73.100 ;
        RECT 59.000 70.800 59.400 71.900 ;
        RECT 60.600 70.800 61.000 72.100 ;
        RECT 62.200 70.800 62.600 72.100 ;
        RECT 64.300 70.800 64.700 73.100 ;
        RECT 67.000 70.800 67.400 72.700 ;
        RECT 70.200 70.800 70.600 74.100 ;
        RECT 74.200 70.800 74.600 72.100 ;
        RECT 77.400 70.800 77.800 74.100 ;
        RECT 78.500 70.800 78.900 73.100 ;
        RECT 80.600 70.800 81.000 72.100 ;
        RECT 82.200 70.800 82.600 72.100 ;
        RECT 83.800 70.800 84.200 71.900 ;
        RECT 88.600 70.800 89.000 73.100 ;
        RECT 91.000 70.800 91.400 73.100 ;
        RECT 93.400 70.800 93.800 73.100 ;
        RECT 95.800 70.800 96.200 73.100 ;
        RECT 0.200 70.200 98.200 70.800 ;
        RECT 3.800 69.100 4.200 70.200 ;
        RECT 5.400 68.900 5.800 70.200 ;
        RECT 8.600 67.900 9.000 70.200 ;
        RECT 9.400 68.900 9.800 70.200 ;
        RECT 11.000 68.900 11.400 70.200 ;
        RECT 14.200 66.900 14.600 70.200 ;
        RECT 16.600 67.900 17.000 70.200 ;
        RECT 19.000 67.900 19.400 70.200 ;
        RECT 19.800 68.900 20.200 70.200 ;
        RECT 21.400 68.900 21.800 70.200 ;
        RECT 22.200 68.900 22.600 70.200 ;
        RECT 23.800 68.900 24.200 70.200 ;
        RECT 24.600 68.900 25.000 70.200 ;
        RECT 26.200 68.900 26.600 70.200 ;
        RECT 28.600 68.900 29.000 70.200 ;
        RECT 30.200 68.900 30.600 70.200 ;
        RECT 31.000 68.900 31.400 70.200 ;
        RECT 32.600 68.900 33.000 70.200 ;
        RECT 33.400 68.900 33.800 70.200 ;
        RECT 35.000 68.900 35.400 70.200 ;
        RECT 35.800 68.900 36.200 70.200 ;
        RECT 37.400 68.900 37.800 70.200 ;
        RECT 38.200 68.900 38.600 70.200 ;
        RECT 39.800 68.900 40.200 70.200 ;
        RECT 40.600 68.900 41.000 70.200 ;
        RECT 42.200 68.900 42.600 70.200 ;
        RECT 43.000 67.900 43.400 70.200 ;
        RECT 44.600 67.900 45.000 70.200 ;
        RECT 47.600 67.900 48.000 70.200 ;
        RECT 50.200 68.300 50.600 70.200 ;
        RECT 51.800 67.900 52.200 70.200 ;
        RECT 53.400 68.900 53.800 70.200 ;
        RECT 55.500 67.900 55.900 70.200 ;
        RECT 58.200 68.300 58.600 70.200 ;
        RECT 60.600 68.300 61.000 70.200 ;
        RECT 63.800 68.900 64.200 70.200 ;
        RECT 65.400 68.900 65.800 70.200 ;
        RECT 66.200 67.900 66.600 70.200 ;
        RECT 69.400 66.900 69.800 70.200 ;
        RECT 72.600 67.900 73.000 70.200 ;
        RECT 75.800 68.300 76.200 70.200 ;
        RECT 78.200 68.900 78.600 70.200 ;
        RECT 79.800 68.900 80.200 70.200 ;
        RECT 80.600 68.900 81.000 70.200 ;
        RECT 82.200 68.900 82.600 70.200 ;
        RECT 85.400 66.900 85.800 70.200 ;
        RECT 86.200 68.900 86.600 70.200 ;
        RECT 88.300 67.900 88.700 70.200 ;
        RECT 89.400 68.900 89.800 70.200 ;
        RECT 91.500 67.900 91.900 70.200 ;
        RECT 93.400 68.900 93.800 70.200 ;
        RECT 95.800 67.900 96.200 70.200 ;
        RECT 0.600 50.800 1.000 53.100 ;
        RECT 3.000 50.800 3.400 54.100 ;
        RECT 7.500 50.800 7.900 53.000 ;
        RECT 11.800 50.800 12.200 52.700 ;
        RECT 13.400 50.800 13.800 53.100 ;
        RECT 15.800 50.800 16.200 53.100 ;
        RECT 18.200 50.800 18.600 52.700 ;
        RECT 20.600 50.800 21.000 54.100 ;
        RECT 25.400 50.800 25.800 52.700 ;
        RECT 28.600 50.800 29.000 52.100 ;
        RECT 30.200 50.800 30.600 52.100 ;
        RECT 32.600 50.800 33.000 53.100 ;
        RECT 33.400 50.800 33.800 52.100 ;
        RECT 35.200 50.800 35.600 53.100 ;
        RECT 38.200 50.800 38.600 53.100 ;
        RECT 40.600 50.800 41.000 52.700 ;
        RECT 42.200 50.800 42.600 52.100 ;
        RECT 43.800 50.800 44.200 52.100 ;
        RECT 46.200 50.800 46.600 52.700 ;
        RECT 47.800 50.800 48.200 52.100 ;
        RECT 51.000 50.800 51.400 53.100 ;
        RECT 53.400 50.800 53.800 52.700 ;
        RECT 56.600 50.800 57.000 52.700 ;
        RECT 58.200 50.800 58.600 52.100 ;
        RECT 59.800 50.800 60.200 52.100 ;
        RECT 63.000 50.800 63.400 52.700 ;
        RECT 65.400 50.800 65.800 52.100 ;
        RECT 66.200 50.800 66.600 52.100 ;
        RECT 67.800 50.800 68.200 52.100 ;
        RECT 70.200 50.800 70.600 52.100 ;
        RECT 71.800 50.800 72.200 52.100 ;
        RECT 72.600 50.800 73.000 54.100 ;
        RECT 75.800 50.800 76.200 52.100 ;
        RECT 77.400 50.800 77.800 52.100 ;
        RECT 78.200 50.800 78.600 52.100 ;
        RECT 79.800 50.800 80.200 52.100 ;
        RECT 82.200 50.800 82.600 52.700 ;
        RECT 83.800 50.800 84.200 52.100 ;
        RECT 85.400 50.800 85.800 52.100 ;
        RECT 87.800 50.800 88.200 52.700 ;
        RECT 90.200 50.800 90.600 52.100 ;
        RECT 91.800 50.800 92.200 53.100 ;
        RECT 93.400 50.800 93.800 53.100 ;
        RECT 95.800 50.800 96.200 52.700 ;
        RECT 0.200 50.200 98.200 50.800 ;
        RECT 0.600 47.900 1.000 50.200 ;
        RECT 2.200 47.900 2.600 50.200 ;
        RECT 5.400 48.300 5.800 50.200 ;
        RECT 9.100 48.000 9.500 50.200 ;
        RECT 11.000 48.900 11.400 50.200 ;
        RECT 12.600 48.900 13.000 50.200 ;
        RECT 13.400 48.900 13.800 50.200 ;
        RECT 15.500 47.900 15.900 50.200 ;
        RECT 17.400 48.100 17.800 50.200 ;
        RECT 19.000 48.900 19.400 50.200 ;
        RECT 20.600 48.300 21.000 50.200 ;
        RECT 23.000 46.900 23.400 50.200 ;
        RECT 27.800 47.900 28.200 50.200 ;
        RECT 31.800 47.900 32.200 50.200 ;
        RECT 32.600 47.900 33.000 50.200 ;
        RECT 35.600 47.900 36.000 50.200 ;
        RECT 36.600 47.900 37.000 50.200 ;
        RECT 39.000 47.900 39.400 50.200 ;
        RECT 42.000 47.900 42.400 50.200 ;
        RECT 44.600 48.300 45.000 50.200 ;
        RECT 46.200 48.900 46.600 50.200 ;
        RECT 47.800 48.900 48.200 50.200 ;
        RECT 48.600 47.900 49.000 50.200 ;
        RECT 51.000 47.900 51.400 50.200 ;
        RECT 53.400 48.300 53.800 50.200 ;
        RECT 55.000 48.900 55.400 50.200 ;
        RECT 57.100 47.900 57.500 50.200 ;
        RECT 58.200 46.900 58.600 50.200 ;
        RECT 62.200 48.300 62.600 50.200 ;
        RECT 65.400 48.300 65.800 50.200 ;
        RECT 69.700 47.900 70.100 50.200 ;
        RECT 71.800 48.900 72.200 50.200 ;
        RECT 72.600 46.900 73.000 50.200 ;
        RECT 75.800 47.900 76.200 50.200 ;
        RECT 78.200 48.300 78.600 50.200 ;
        RECT 80.900 47.900 81.300 50.200 ;
        RECT 83.000 48.900 83.400 50.200 ;
        RECT 83.800 48.900 84.200 50.200 ;
        RECT 85.400 48.900 85.800 50.200 ;
        RECT 89.400 49.100 89.800 50.200 ;
        RECT 91.000 48.900 91.400 50.200 ;
        RECT 93.400 47.900 93.800 50.200 ;
        RECT 96.300 48.000 96.700 50.200 ;
        RECT 1.400 30.800 1.800 32.700 ;
        RECT 4.000 30.800 4.400 33.100 ;
        RECT 7.000 30.800 7.400 33.100 ;
        RECT 7.800 30.800 8.200 33.100 ;
        RECT 10.200 30.800 10.600 32.700 ;
        RECT 12.600 30.800 13.000 32.100 ;
        RECT 14.200 30.800 14.600 32.100 ;
        RECT 15.000 30.800 15.400 32.100 ;
        RECT 16.600 30.800 17.000 32.900 ;
        RECT 18.500 30.800 18.900 33.100 ;
        RECT 20.600 30.800 21.000 32.100 ;
        RECT 21.700 30.800 22.100 33.100 ;
        RECT 23.800 30.800 24.200 32.100 ;
        RECT 24.600 30.800 25.000 32.100 ;
        RECT 26.200 30.800 26.600 32.100 ;
        RECT 29.400 30.800 29.800 32.700 ;
        RECT 33.400 30.800 33.800 33.100 ;
        RECT 34.500 30.800 34.900 33.100 ;
        RECT 36.600 30.800 37.000 32.100 ;
        RECT 38.200 30.800 38.600 32.700 ;
        RECT 41.400 30.800 41.800 32.100 ;
        RECT 42.200 30.800 42.600 32.100 ;
        RECT 43.800 30.800 44.200 32.100 ;
        RECT 45.400 30.800 45.800 32.700 ;
        RECT 47.800 30.800 48.200 32.100 ;
        RECT 49.400 30.800 49.800 32.100 ;
        RECT 50.400 30.800 50.800 33.100 ;
        RECT 53.400 30.800 53.800 33.100 ;
        RECT 55.800 30.800 56.200 32.700 ;
        RECT 58.200 30.800 58.600 32.100 ;
        RECT 62.200 30.800 62.600 31.900 ;
        RECT 63.800 30.800 64.200 32.100 ;
        RECT 66.200 30.800 66.600 32.700 ;
        RECT 71.800 30.800 72.200 32.700 ;
        RECT 75.000 30.800 75.400 33.100 ;
        RECT 76.600 30.800 77.000 32.700 ;
        RECT 79.000 30.800 79.400 32.100 ;
        RECT 82.200 30.800 82.600 32.700 ;
        RECT 85.400 30.800 85.800 32.700 ;
        RECT 87.800 30.800 88.200 33.100 ;
        RECT 89.400 30.800 89.800 32.700 ;
        RECT 91.800 30.800 92.200 32.100 ;
        RECT 95.000 30.800 95.400 33.100 ;
        RECT 0.200 30.200 98.200 30.800 ;
        RECT 1.400 27.900 1.800 30.200 ;
        RECT 4.600 27.900 5.000 30.200 ;
        RECT 7.800 26.900 8.200 30.200 ;
        RECT 10.200 28.300 10.600 30.200 ;
        RECT 15.000 29.100 15.400 30.200 ;
        RECT 16.600 28.900 17.000 30.200 ;
        RECT 19.800 28.300 20.200 30.200 ;
        RECT 23.000 28.300 23.400 30.200 ;
        RECT 24.600 28.900 25.000 30.200 ;
        RECT 26.200 28.100 26.600 30.200 ;
        RECT 29.400 28.900 29.800 30.200 ;
        RECT 31.000 28.900 31.400 30.200 ;
        RECT 31.800 26.900 32.200 30.200 ;
        RECT 35.800 28.300 36.200 30.200 ;
        RECT 39.000 28.900 39.400 30.200 ;
        RECT 39.800 28.900 40.200 30.200 ;
        RECT 41.400 28.900 41.800 30.200 ;
        RECT 43.000 28.300 43.400 30.200 ;
        RECT 46.200 28.900 46.600 30.200 ;
        RECT 47.200 27.900 47.600 30.200 ;
        RECT 50.200 27.900 50.600 30.200 ;
        RECT 51.000 28.900 51.400 30.200 ;
        RECT 52.600 27.900 53.000 30.200 ;
        RECT 55.600 27.900 56.000 30.200 ;
        RECT 56.900 27.900 57.300 30.200 ;
        RECT 59.000 28.900 59.400 30.200 ;
        RECT 60.100 27.900 60.500 30.200 ;
        RECT 62.200 28.900 62.600 30.200 ;
        RECT 63.800 28.300 64.200 30.200 ;
        RECT 66.200 28.900 66.600 30.200 ;
        RECT 67.800 28.900 68.200 30.200 ;
        RECT 71.800 28.300 72.200 30.200 ;
        RECT 75.000 27.900 75.400 30.200 ;
        RECT 77.400 28.300 77.800 30.200 ;
        RECT 79.000 28.900 79.400 30.200 ;
        RECT 80.600 28.900 81.000 30.200 ;
        RECT 81.700 27.900 82.100 30.200 ;
        RECT 83.800 28.900 84.200 30.200 ;
        RECT 86.200 28.300 86.600 30.200 ;
        RECT 88.600 27.900 89.000 30.200 ;
        RECT 91.000 27.900 91.400 30.200 ;
        RECT 91.800 28.900 92.200 30.200 ;
        RECT 93.400 28.900 93.800 30.200 ;
        RECT 95.800 28.300 96.200 30.200 ;
        RECT 3.800 10.800 4.200 11.900 ;
        RECT 5.400 10.800 5.800 12.100 ;
        RECT 7.800 10.800 8.200 12.700 ;
        RECT 12.600 10.800 13.000 14.100 ;
        RECT 13.400 10.800 13.800 13.100 ;
        RECT 17.400 10.800 17.800 13.100 ;
        RECT 18.500 10.800 18.900 13.100 ;
        RECT 20.600 10.800 21.000 12.100 ;
        RECT 23.000 10.800 23.400 12.700 ;
        RECT 24.600 10.800 25.000 13.100 ;
        RECT 28.600 10.800 29.000 13.100 ;
        RECT 31.000 10.800 31.400 14.100 ;
        RECT 35.000 10.800 35.400 12.700 ;
        RECT 37.400 10.800 37.800 12.100 ;
        RECT 39.000 10.800 39.400 12.100 ;
        RECT 39.800 10.800 40.200 12.100 ;
        RECT 41.900 10.800 42.300 13.100 ;
        RECT 43.300 10.800 43.700 13.100 ;
        RECT 45.400 10.800 45.800 12.100 ;
        RECT 48.600 10.800 49.000 14.100 ;
        RECT 49.400 10.800 49.800 13.100 ;
        RECT 52.400 10.800 52.800 13.100 ;
        RECT 54.200 10.800 54.600 12.700 ;
        RECT 57.400 10.800 57.800 12.100 ;
        RECT 59.000 10.800 59.400 11.900 ;
        RECT 63.800 10.800 64.200 12.700 ;
        RECT 67.800 10.800 68.200 12.700 ;
        RECT 71.000 10.800 71.400 13.100 ;
        RECT 72.600 10.800 73.000 12.100 ;
        RECT 74.200 10.800 74.600 12.100 ;
        RECT 75.800 10.800 76.200 13.100 ;
        RECT 76.900 10.800 77.300 13.100 ;
        RECT 79.000 10.800 79.400 12.100 ;
        RECT 81.400 10.800 81.800 12.700 ;
        RECT 83.800 10.800 84.200 12.700 ;
        RECT 86.200 10.800 86.600 12.100 ;
        RECT 88.300 10.800 88.700 13.100 ;
        RECT 89.400 10.800 89.800 14.100 ;
        RECT 92.600 10.800 93.000 12.100 ;
        RECT 94.700 10.800 95.100 13.100 ;
        RECT 0.200 10.200 98.200 10.800 ;
        RECT 1.400 8.200 1.900 10.200 ;
        RECT 4.500 9.900 4.900 10.200 ;
        RECT 4.500 8.200 5.000 9.900 ;
        RECT 7.500 8.000 7.900 10.200 ;
        RECT 9.400 8.900 9.800 10.200 ;
        RECT 11.000 8.100 11.400 10.200 ;
        RECT 14.200 7.900 14.600 10.200 ;
        RECT 15.200 7.900 15.600 10.200 ;
        RECT 18.200 7.900 18.600 10.200 ;
        RECT 20.600 7.900 21.000 10.200 ;
        RECT 21.400 8.900 21.800 10.200 ;
        RECT 23.000 8.900 23.400 10.200 ;
        RECT 24.600 8.300 25.000 10.200 ;
        RECT 29.400 8.900 29.800 10.200 ;
        RECT 31.000 8.900 31.400 10.200 ;
        RECT 32.600 8.300 33.000 10.200 ;
        RECT 36.600 7.900 37.000 10.200 ;
        RECT 38.200 8.100 38.600 10.200 ;
        RECT 39.800 8.900 40.200 10.200 ;
        RECT 40.800 7.900 41.200 10.200 ;
        RECT 43.800 7.900 44.200 10.200 ;
        RECT 45.700 8.000 46.100 10.200 ;
        RECT 48.700 9.900 49.100 10.200 ;
        RECT 48.600 8.200 49.100 9.900 ;
        RECT 51.700 8.200 52.200 10.200 ;
        RECT 54.200 7.900 54.600 10.200 ;
        RECT 56.600 7.900 57.000 10.200 ;
        RECT 59.000 8.200 59.500 10.200 ;
        RECT 62.100 9.900 62.500 10.200 ;
        RECT 62.100 8.200 62.600 9.900 ;
        RECT 63.800 7.900 64.200 10.200 ;
        RECT 66.800 7.900 67.200 10.200 ;
        RECT 71.000 7.900 71.400 10.200 ;
        RECT 71.800 7.900 72.200 10.200 ;
        RECT 73.400 7.900 73.800 10.200 ;
        RECT 75.800 8.900 76.200 10.200 ;
        RECT 78.200 8.300 78.600 10.200 ;
        RECT 81.400 7.900 81.800 10.200 ;
        RECT 82.200 7.900 82.600 10.200 ;
        RECT 84.600 8.900 85.000 10.200 ;
        RECT 86.200 8.900 86.600 10.200 ;
        RECT 87.800 7.900 88.200 10.200 ;
        RECT 90.200 8.900 90.600 10.200 ;
        RECT 91.800 8.200 92.300 10.200 ;
        RECT 94.900 9.900 95.300 10.200 ;
        RECT 94.900 8.200 95.400 9.900 ;
      LAYER via1 ;
        RECT 68.200 70.300 68.600 70.700 ;
        RECT 68.900 70.300 69.300 70.700 ;
        RECT 68.200 50.300 68.600 50.700 ;
        RECT 68.900 50.300 69.300 50.700 ;
        RECT 68.200 30.300 68.600 30.700 ;
        RECT 68.900 30.300 69.300 30.700 ;
        RECT 68.200 10.300 68.600 10.700 ;
        RECT 68.900 10.300 69.300 10.700 ;
      LAYER metal2 ;
        RECT 68.000 70.300 69.600 70.700 ;
        RECT 68.000 50.300 69.600 50.700 ;
        RECT 68.000 30.300 69.600 30.700 ;
        RECT 68.000 10.300 69.600 10.700 ;
      LAYER via2 ;
        RECT 68.200 70.300 68.600 70.700 ;
        RECT 68.900 70.300 69.300 70.700 ;
        RECT 68.200 50.300 68.600 50.700 ;
        RECT 68.900 50.300 69.300 50.700 ;
        RECT 68.200 30.300 68.600 30.700 ;
        RECT 68.900 30.300 69.300 30.700 ;
        RECT 68.200 10.300 68.600 10.700 ;
        RECT 68.900 10.300 69.300 10.700 ;
      LAYER metal3 ;
        RECT 68.000 70.300 69.600 70.700 ;
        RECT 68.000 50.300 69.600 50.700 ;
        RECT 68.000 30.300 69.600 30.700 ;
        RECT 68.000 10.300 69.600 10.700 ;
      LAYER via3 ;
        RECT 68.200 70.300 68.600 70.700 ;
        RECT 69.000 70.300 69.400 70.700 ;
        RECT 68.200 50.300 68.600 50.700 ;
        RECT 69.000 50.300 69.400 50.700 ;
        RECT 68.200 30.300 68.600 30.700 ;
        RECT 69.000 30.300 69.400 30.700 ;
        RECT 68.200 10.300 68.600 10.700 ;
        RECT 69.000 10.300 69.400 10.700 ;
      LAYER metal4 ;
        RECT 68.000 70.300 69.600 70.700 ;
        RECT 68.000 50.300 69.600 50.700 ;
        RECT 68.000 30.300 69.600 30.700 ;
        RECT 68.000 10.300 69.600 10.700 ;
      LAYER via4 ;
        RECT 68.200 70.300 68.600 70.700 ;
        RECT 68.900 70.300 69.300 70.700 ;
        RECT 68.200 50.300 68.600 50.700 ;
        RECT 68.900 50.300 69.300 50.700 ;
        RECT 68.200 30.300 68.600 30.700 ;
        RECT 68.900 30.300 69.300 30.700 ;
        RECT 68.200 10.300 68.600 10.700 ;
        RECT 68.900 10.300 69.300 10.700 ;
      LAYER metal5 ;
        RECT 68.000 70.200 69.600 70.700 ;
        RECT 68.000 50.200 69.600 50.700 ;
        RECT 68.000 30.200 69.600 30.700 ;
        RECT 68.000 10.200 69.600 10.700 ;
      LAYER via5 ;
        RECT 69.000 70.200 69.500 70.700 ;
        RECT 69.000 50.200 69.500 50.700 ;
        RECT 69.000 30.200 69.500 30.700 ;
        RECT 69.000 10.200 69.500 10.700 ;
      LAYER metal6 ;
        RECT 68.000 -3.000 69.600 83.000 ;
    END
  END gnd
  PIN A[0]
    PORT
      LAYER metal1 ;
        RECT 13.400 54.800 13.800 55.200 ;
        RECT 0.600 53.400 1.000 54.200 ;
        RECT 6.200 53.800 6.600 54.600 ;
        RECT 13.400 54.200 13.700 54.800 ;
        RECT 12.600 54.100 13.000 54.200 ;
        RECT 13.400 54.100 13.800 54.200 ;
        RECT 12.200 53.800 13.800 54.100 ;
        RECT 12.200 53.600 12.600 53.800 ;
        RECT 13.400 53.400 13.800 53.800 ;
        RECT 15.800 53.400 16.200 54.200 ;
      LAYER via1 ;
        RECT 0.600 53.800 1.000 54.200 ;
        RECT 15.800 53.800 16.200 54.200 ;
      LAYER metal2 ;
        RECT 0.600 56.800 1.000 57.200 ;
        RECT 0.600 54.200 0.900 56.800 ;
        RECT 13.400 54.800 13.800 55.200 ;
        RECT 13.400 54.200 13.700 54.800 ;
        RECT 0.600 54.100 1.000 54.200 ;
        RECT 1.400 54.100 1.800 54.200 ;
        RECT 0.600 53.800 1.800 54.100 ;
        RECT 6.200 54.100 6.600 54.200 ;
        RECT 7.000 54.100 7.400 54.200 ;
        RECT 6.200 53.800 7.400 54.100 ;
        RECT 13.400 53.800 13.800 54.200 ;
        RECT 15.000 54.100 15.400 54.200 ;
        RECT 15.800 54.100 16.200 54.200 ;
        RECT 15.000 53.800 16.200 54.100 ;
      LAYER via2 ;
        RECT 1.400 53.800 1.800 54.200 ;
        RECT 7.000 53.800 7.400 54.200 ;
      LAYER metal3 ;
        RECT -2.600 57.100 -2.200 57.200 ;
        RECT 0.600 57.100 1.000 57.200 ;
        RECT -2.600 56.800 1.000 57.100 ;
        RECT 1.400 54.100 1.800 54.200 ;
        RECT 7.000 54.100 7.400 54.200 ;
        RECT 13.400 54.100 13.800 54.200 ;
        RECT 15.000 54.100 15.400 54.200 ;
        RECT 1.400 53.800 15.400 54.100 ;
    END
  END A[0]
  PIN A[1]
    PORT
      LAYER metal1 ;
        RECT 12.600 47.800 13.000 48.600 ;
        RECT 19.000 47.800 19.400 48.600 ;
        RECT 0.600 46.800 1.000 47.600 ;
        RECT 5.000 47.200 5.400 47.400 ;
        RECT 4.600 46.900 5.400 47.200 ;
        RECT 4.600 46.800 5.000 46.900 ;
        RECT 7.800 46.400 8.200 47.200 ;
        RECT 27.800 46.800 28.200 47.600 ;
        RECT 41.400 46.400 41.800 47.200 ;
      LAYER via1 ;
        RECT 7.800 46.800 8.200 47.200 ;
        RECT 41.400 46.800 41.800 47.200 ;
      LAYER metal2 ;
        RECT 0.600 47.800 1.000 48.200 ;
        RECT 4.600 47.800 5.000 48.200 ;
        RECT 12.600 47.800 13.000 48.200 ;
        RECT 19.000 47.800 19.400 48.200 ;
        RECT 0.600 47.200 0.900 47.800 ;
        RECT 4.600 47.200 4.900 47.800 ;
        RECT 12.600 47.200 12.900 47.800 ;
        RECT 19.000 47.200 19.300 47.800 ;
        RECT 0.600 46.800 1.000 47.200 ;
        RECT 4.600 46.800 5.000 47.200 ;
        RECT 7.800 47.100 8.200 47.200 ;
        RECT 8.600 47.100 9.000 47.200 ;
        RECT 7.800 46.800 9.000 47.100 ;
        RECT 12.600 46.800 13.000 47.200 ;
        RECT 19.000 46.800 19.400 47.200 ;
        RECT 27.000 47.100 27.400 47.200 ;
        RECT 27.800 47.100 28.200 47.200 ;
        RECT 27.000 46.800 28.200 47.100 ;
        RECT 40.600 47.100 41.000 47.200 ;
        RECT 41.400 47.100 41.800 47.200 ;
        RECT 40.600 46.800 41.800 47.100 ;
      LAYER via2 ;
        RECT 8.600 46.800 9.000 47.200 ;
      LAYER metal3 ;
        RECT 0.600 47.800 1.000 48.200 ;
        RECT 4.600 47.800 5.000 48.200 ;
        RECT -2.600 47.100 -2.200 47.200 ;
        RECT 0.600 47.100 0.900 47.800 ;
        RECT 4.600 47.100 4.900 47.800 ;
        RECT 8.600 47.100 9.000 47.200 ;
        RECT 12.600 47.100 13.000 47.200 ;
        RECT 19.000 47.100 19.400 47.200 ;
        RECT 27.000 47.100 27.400 47.200 ;
        RECT 40.600 47.100 41.000 47.200 ;
        RECT -2.600 46.800 41.000 47.100 ;
    END
  END A[1]
  PIN A[2]
    PORT
      LAYER metal1 ;
        RECT 19.000 66.800 19.400 67.600 ;
        RECT 7.800 33.400 8.200 34.200 ;
        RECT 26.200 16.100 26.600 16.600 ;
        RECT 27.000 16.100 27.400 16.200 ;
        RECT 26.200 15.800 27.400 16.100 ;
        RECT 7.000 15.100 7.400 15.200 ;
        RECT 7.800 15.100 8.200 15.200 ;
        RECT 7.000 14.800 8.200 15.100 ;
        RECT 49.400 14.800 49.800 15.600 ;
        RECT 7.800 14.400 8.200 14.800 ;
        RECT 0.600 6.800 1.400 7.200 ;
        RECT 7.200 6.900 7.600 7.000 ;
        RECT 7.100 6.600 7.600 6.900 ;
        RECT 10.200 6.800 10.700 7.200 ;
        RECT 7.100 6.200 7.400 6.600 ;
        RECT 10.400 6.400 10.800 6.800 ;
        RECT 7.000 5.800 7.400 6.200 ;
        RECT 21.400 5.400 21.800 6.200 ;
      LAYER via1 ;
        RECT 7.800 33.800 8.200 34.200 ;
        RECT 27.000 15.800 27.400 16.200 ;
        RECT 21.400 5.800 21.800 6.200 ;
      LAYER metal2 ;
        RECT 18.200 67.100 18.600 67.200 ;
        RECT 19.000 67.100 19.400 67.200 ;
        RECT 18.200 66.800 19.400 67.100 ;
        RECT 7.800 33.800 8.200 34.200 ;
        RECT 7.800 21.100 8.100 33.800 ;
        RECT 7.000 20.800 8.100 21.100 ;
        RECT 7.000 15.200 7.300 20.800 ;
        RECT 27.000 17.800 27.400 18.200 ;
        RECT 49.400 17.800 49.800 18.200 ;
        RECT 27.000 16.200 27.300 17.800 ;
        RECT 27.000 15.800 27.400 16.200 ;
        RECT 7.000 14.800 7.400 15.200 ;
        RECT 7.000 9.200 7.300 14.800 ;
        RECT 27.000 12.200 27.300 15.800 ;
        RECT 49.400 15.200 49.700 17.800 ;
        RECT 49.400 14.800 49.800 15.200 ;
        RECT 21.400 11.800 21.800 12.200 ;
        RECT 27.000 11.800 27.400 12.200 ;
        RECT 0.600 8.800 1.000 9.200 ;
        RECT 7.000 8.800 7.400 9.200 ;
        RECT 10.200 8.800 10.600 9.200 ;
        RECT 0.600 7.200 0.900 8.800 ;
        RECT 0.600 6.800 1.000 7.200 ;
        RECT 7.000 6.200 7.300 8.800 ;
        RECT 10.200 7.200 10.500 8.800 ;
        RECT 21.400 7.200 21.700 11.800 ;
        RECT 10.200 6.800 10.600 7.200 ;
        RECT 21.400 6.800 21.800 7.200 ;
        RECT 21.400 6.200 21.700 6.800 ;
        RECT 7.000 5.800 7.400 6.200 ;
        RECT 21.400 5.800 21.800 6.200 ;
      LAYER metal3 ;
        RECT 18.200 67.100 18.600 67.200 ;
        RECT 19.000 67.100 19.400 67.200 ;
        RECT 18.200 66.800 19.400 67.100 ;
        RECT 7.800 34.100 8.200 34.200 ;
        RECT 19.000 34.100 19.400 34.200 ;
        RECT 7.800 33.800 19.400 34.100 ;
        RECT 27.000 18.100 27.400 18.200 ;
        RECT 49.400 18.100 49.800 18.200 ;
        RECT 27.000 17.800 49.800 18.100 ;
        RECT 21.400 12.100 21.800 12.200 ;
        RECT 27.000 12.100 27.400 12.200 ;
        RECT 21.400 11.800 27.400 12.100 ;
        RECT -2.600 9.100 -2.200 9.200 ;
        RECT 0.600 9.100 1.000 9.200 ;
        RECT 7.000 9.100 7.400 9.200 ;
        RECT 10.200 9.100 10.600 9.200 ;
        RECT -2.600 8.800 10.600 9.100 ;
        RECT 10.200 7.100 10.600 7.200 ;
        RECT 21.400 7.100 21.800 7.200 ;
        RECT 10.200 6.800 21.800 7.100 ;
      LAYER via3 ;
        RECT 19.000 66.800 19.400 67.200 ;
        RECT 19.000 33.800 19.400 34.200 ;
      LAYER metal4 ;
        RECT 19.000 66.800 19.400 67.200 ;
        RECT 19.000 34.200 19.300 66.800 ;
        RECT 19.000 33.800 19.400 34.200 ;
    END
  END A[2]
  PIN A[3]
    PORT
      LAYER metal1 ;
        RECT 46.200 27.800 46.600 28.600 ;
        RECT 52.600 25.400 53.000 26.200 ;
        RECT 17.400 14.100 17.800 14.200 ;
        RECT 18.200 14.100 18.600 14.200 ;
        RECT 17.400 13.800 18.600 14.100 ;
        RECT 17.400 13.400 17.800 13.800 ;
        RECT 38.900 6.800 39.400 7.200 ;
        RECT 38.800 6.400 39.200 6.800 ;
        RECT 46.000 6.600 46.600 7.000 ;
        RECT 52.200 6.800 53.000 7.200 ;
        RECT 46.200 6.200 46.500 6.600 ;
        RECT 29.400 5.400 29.800 6.200 ;
        RECT 46.200 5.800 46.600 6.200 ;
        RECT 35.000 4.400 35.400 5.200 ;
      LAYER via1 ;
        RECT 52.600 25.800 53.000 26.200 ;
        RECT 18.200 13.800 18.600 14.200 ;
        RECT 39.000 6.800 39.400 7.200 ;
        RECT 46.200 6.600 46.600 7.000 ;
        RECT 52.600 6.800 53.000 7.200 ;
        RECT 29.400 5.800 29.800 6.200 ;
        RECT 35.000 4.800 35.400 5.200 ;
      LAYER metal2 ;
        RECT 46.200 27.800 46.600 28.200 ;
        RECT 46.200 27.200 46.500 27.800 ;
        RECT 46.200 26.800 46.600 27.200 ;
        RECT 52.600 26.800 53.000 27.200 ;
        RECT 18.200 13.800 18.600 14.200 ;
        RECT 18.200 8.200 18.500 13.800 ;
        RECT 46.200 8.200 46.500 26.800 ;
        RECT 52.600 26.200 52.900 26.800 ;
        RECT 52.600 25.800 53.000 26.200 ;
        RECT 18.200 7.800 18.600 8.200 ;
        RECT 29.400 7.800 29.800 8.200 ;
        RECT 35.000 7.800 35.400 8.200 ;
        RECT 39.000 7.800 39.400 8.200 ;
        RECT 46.200 7.800 46.600 8.200 ;
        RECT 52.600 7.800 53.000 8.200 ;
        RECT 29.400 6.200 29.700 7.800 ;
        RECT 29.400 5.800 29.800 6.200 ;
        RECT 35.000 5.200 35.300 7.800 ;
        RECT 39.000 7.200 39.300 7.800 ;
        RECT 39.000 6.800 39.400 7.200 ;
        RECT 46.200 7.000 46.500 7.800 ;
        RECT 52.600 7.200 52.900 7.800 ;
        RECT 46.200 6.600 46.600 7.000 ;
        RECT 52.600 6.800 53.000 7.200 ;
        RECT 35.000 4.800 35.400 5.200 ;
        RECT 35.000 2.200 35.300 4.800 ;
        RECT 33.400 1.800 33.800 2.200 ;
        RECT 35.000 1.800 35.400 2.200 ;
        RECT 33.400 -1.800 33.700 1.800 ;
        RECT 33.400 -2.200 33.800 -1.800 ;
      LAYER metal3 ;
        RECT 46.200 27.100 46.600 27.200 ;
        RECT 52.600 27.100 53.000 27.200 ;
        RECT 46.200 26.800 53.000 27.100 ;
        RECT 18.200 8.100 18.600 8.200 ;
        RECT 29.400 8.100 29.800 8.200 ;
        RECT 35.000 8.100 35.400 8.200 ;
        RECT 39.000 8.100 39.400 8.200 ;
        RECT 46.200 8.100 46.600 8.200 ;
        RECT 52.600 8.100 53.000 8.200 ;
        RECT 18.200 7.800 53.000 8.100 ;
        RECT 33.400 2.100 33.800 2.200 ;
        RECT 35.000 2.100 35.400 2.200 ;
        RECT 33.400 1.800 35.400 2.100 ;
    END
  END A[3]
  PIN A[4]
    PORT
      LAYER metal1 ;
        RECT 51.800 14.100 52.200 14.600 ;
        RECT 52.600 14.100 53.000 14.200 ;
        RECT 51.800 13.800 53.000 14.100 ;
        RECT 58.200 6.800 59.000 7.200 ;
        RECT 81.400 7.100 81.800 7.600 ;
        RECT 82.200 7.100 82.600 7.600 ;
        RECT 81.400 6.800 82.600 7.100 ;
        RECT 75.000 4.400 75.400 5.200 ;
      LAYER via1 ;
        RECT 52.600 13.800 53.000 14.200 ;
        RECT 75.000 4.800 75.400 5.200 ;
      LAYER metal2 ;
        RECT 52.600 13.800 53.000 14.200 ;
        RECT 52.600 9.200 52.900 13.800 ;
        RECT 52.600 8.800 53.000 9.200 ;
        RECT 58.200 8.800 58.600 9.200 ;
        RECT 58.200 7.200 58.500 8.800 ;
        RECT 58.200 6.800 58.600 7.200 ;
        RECT 81.400 6.800 81.800 7.200 ;
        RECT 58.200 1.200 58.500 6.800 ;
        RECT 75.000 4.800 75.400 5.200 ;
        RECT 75.000 1.200 75.300 4.800 ;
        RECT 81.400 1.200 81.700 6.800 ;
        RECT 58.200 0.800 58.600 1.200 ;
        RECT 73.400 0.800 73.800 1.200 ;
        RECT 75.000 0.800 75.400 1.200 ;
        RECT 81.400 0.800 81.800 1.200 ;
        RECT 73.400 -1.800 73.700 0.800 ;
        RECT 73.400 -2.200 73.800 -1.800 ;
      LAYER metal3 ;
        RECT 52.600 9.100 53.000 9.200 ;
        RECT 58.200 9.100 58.600 9.200 ;
        RECT 52.600 8.800 58.600 9.100 ;
        RECT 58.200 1.100 58.600 1.200 ;
        RECT 73.400 1.100 73.800 1.200 ;
        RECT 75.000 1.100 75.400 1.200 ;
        RECT 81.400 1.100 81.800 1.200 ;
        RECT 58.200 0.800 81.800 1.100 ;
    END
  END A[4]
  PIN A[5]
    PORT
      LAYER metal1 ;
        RECT 57.400 46.100 57.800 46.200 ;
        RECT 57.000 45.800 57.800 46.100 ;
        RECT 57.000 45.600 57.400 45.800 ;
        RECT 73.400 35.800 73.800 36.600 ;
        RECT 71.800 35.100 72.200 35.200 ;
        RECT 73.400 35.100 73.700 35.800 ;
        RECT 71.800 34.800 73.700 35.100 ;
        RECT 71.800 34.400 72.200 34.800 ;
        RECT 95.000 33.400 95.400 34.200 ;
        RECT 58.200 32.400 58.600 33.200 ;
        RECT 91.000 6.800 91.800 7.200 ;
      LAYER via1 ;
        RECT 57.400 45.800 57.800 46.200 ;
        RECT 95.000 33.800 95.400 34.200 ;
        RECT 58.200 32.800 58.600 33.200 ;
      LAYER metal2 ;
        RECT 57.400 46.100 57.800 46.200 ;
        RECT 57.400 45.800 58.500 46.100 ;
        RECT 58.200 35.200 58.500 45.800 ;
        RECT 58.200 34.800 58.600 35.200 ;
        RECT 71.000 35.100 71.400 35.200 ;
        RECT 71.800 35.100 72.200 35.200 ;
        RECT 71.000 34.800 72.200 35.100 ;
        RECT 95.000 34.800 95.400 35.200 ;
        RECT 58.200 33.200 58.500 34.800 ;
        RECT 71.800 34.200 72.100 34.800 ;
        RECT 95.000 34.200 95.300 34.800 ;
        RECT 71.800 33.800 72.200 34.200 ;
        RECT 95.000 33.800 95.400 34.200 ;
        RECT 58.200 32.800 58.600 33.200 ;
        RECT 91.000 7.800 91.400 8.200 ;
        RECT 91.000 7.200 91.300 7.800 ;
        RECT 91.000 6.800 91.400 7.200 ;
      LAYER metal3 ;
        RECT 58.200 35.100 58.600 35.200 ;
        RECT 71.000 35.100 71.400 35.200 ;
        RECT 58.200 34.800 71.400 35.100 ;
        RECT 95.000 34.800 95.400 35.200 ;
        RECT 71.800 34.100 72.200 34.200 ;
        RECT 91.000 34.100 91.400 34.200 ;
        RECT 95.000 34.100 95.300 34.800 ;
        RECT 100.600 34.100 101.000 34.200 ;
        RECT 71.800 33.800 101.000 34.100 ;
        RECT 91.000 7.800 91.400 8.200 ;
        RECT 91.000 7.200 91.300 7.800 ;
        RECT 91.000 6.800 91.400 7.200 ;
      LAYER via3 ;
        RECT 91.000 33.800 91.400 34.200 ;
      LAYER metal4 ;
        RECT 91.000 33.800 91.400 34.200 ;
        RECT 91.000 7.200 91.300 33.800 ;
        RECT 91.000 6.800 91.400 7.200 ;
    END
  END A[5]
  PIN A[6]
    PORT
      LAYER metal1 ;
        RECT 79.800 54.800 80.200 55.600 ;
        RECT 91.800 53.400 92.200 54.200 ;
        RECT 51.000 33.800 51.400 34.600 ;
      LAYER via1 ;
        RECT 91.800 53.800 92.200 54.200 ;
      LAYER metal2 ;
        RECT 91.800 57.800 92.200 58.200 ;
        RECT 79.800 54.800 80.200 55.200 ;
        RECT 79.800 52.200 80.100 54.800 ;
        RECT 91.800 54.200 92.100 57.800 ;
        RECT 91.800 53.800 92.200 54.200 ;
        RECT 91.800 52.200 92.100 53.800 ;
        RECT 79.800 51.800 80.200 52.200 ;
        RECT 91.800 51.800 92.200 52.200 ;
        RECT 51.800 50.800 52.200 51.200 ;
        RECT 51.800 46.100 52.100 50.800 ;
        RECT 51.000 45.800 52.100 46.100 ;
        RECT 51.000 34.200 51.300 45.800 ;
        RECT 51.000 33.800 51.400 34.200 ;
      LAYER metal3 ;
        RECT 91.800 58.100 92.200 58.200 ;
        RECT 100.600 58.100 101.000 58.200 ;
        RECT 91.800 57.800 101.000 58.100 ;
        RECT 79.800 52.100 80.200 52.200 ;
        RECT 91.800 52.100 92.200 52.200 ;
        RECT 67.000 51.800 92.200 52.100 ;
        RECT 51.800 51.100 52.200 51.200 ;
        RECT 67.000 51.100 67.300 51.800 ;
        RECT 51.800 50.800 67.300 51.100 ;
    END
  END A[6]
  PIN A[7]
    PORT
      LAYER metal1 ;
        RECT 41.800 75.200 42.200 75.400 ;
        RECT 41.800 74.900 42.600 75.200 ;
        RECT 42.200 74.800 42.600 74.900 ;
        RECT 50.200 74.800 50.600 75.600 ;
        RECT 47.800 73.400 48.200 74.200 ;
        RECT 59.000 73.800 60.200 74.200 ;
      LAYER via1 ;
        RECT 47.800 73.800 48.200 74.200 ;
      LAYER metal2 ;
        RECT 49.400 82.800 49.800 83.200 ;
        RECT 49.400 75.200 49.700 82.800 ;
        RECT 42.200 75.100 42.600 75.200 ;
        RECT 43.000 75.100 43.400 75.200 ;
        RECT 42.200 74.800 43.400 75.100 ;
        RECT 47.800 74.800 48.200 75.200 ;
        RECT 49.400 75.100 49.800 75.200 ;
        RECT 50.200 75.100 50.600 75.200 ;
        RECT 49.400 74.800 50.600 75.100 ;
        RECT 59.000 74.800 59.400 75.200 ;
        RECT 47.800 74.200 48.100 74.800 ;
        RECT 59.000 74.200 59.300 74.800 ;
        RECT 47.800 73.800 48.200 74.200 ;
        RECT 59.000 73.800 59.400 74.200 ;
      LAYER via2 ;
        RECT 43.000 74.800 43.400 75.200 ;
      LAYER metal3 ;
        RECT 43.000 75.100 43.400 75.200 ;
        RECT 47.800 75.100 48.200 75.200 ;
        RECT 49.400 75.100 49.800 75.200 ;
        RECT 59.000 75.100 59.400 75.200 ;
        RECT 43.000 74.800 59.400 75.100 ;
    END
  END A[7]
  PIN B[0]
    PORT
      LAYER metal1 ;
        RECT 15.000 55.800 15.400 56.600 ;
        RECT 7.000 54.800 7.400 55.200 ;
        RECT 7.100 54.400 7.400 54.800 ;
        RECT 7.100 54.100 7.600 54.400 ;
        RECT 7.200 54.000 7.600 54.100 ;
        RECT 32.600 54.100 33.000 54.200 ;
        RECT 32.600 53.800 33.700 54.100 ;
        RECT 32.600 53.400 33.000 53.800 ;
        RECT 33.400 53.200 33.700 53.800 ;
        RECT 33.400 52.400 33.800 53.200 ;
        RECT 35.000 46.400 35.400 47.200 ;
      LAYER via1 ;
        RECT 33.400 52.800 33.800 53.200 ;
        RECT 35.000 46.800 35.400 47.200 ;
      LAYER metal2 ;
        RECT 15.000 55.800 15.400 56.200 ;
        RECT 15.000 55.200 15.300 55.800 ;
        RECT 7.000 55.100 7.400 55.200 ;
        RECT 7.800 55.100 8.200 55.200 ;
        RECT 7.000 54.800 8.200 55.100 ;
        RECT 15.000 54.800 15.400 55.200 ;
        RECT 33.400 54.800 33.800 55.200 ;
        RECT 33.400 53.200 33.700 54.800 ;
        RECT 33.400 53.100 33.800 53.200 ;
        RECT 34.200 53.100 34.600 53.200 ;
        RECT 33.400 52.800 34.600 53.100 ;
        RECT 35.000 52.800 35.400 53.200 ;
        RECT 35.000 47.200 35.300 52.800 ;
        RECT 35.000 46.800 35.400 47.200 ;
      LAYER via2 ;
        RECT 7.800 54.800 8.200 55.200 ;
        RECT 34.200 52.800 34.600 53.200 ;
      LAYER metal3 ;
        RECT -2.600 55.100 -2.200 55.200 ;
        RECT 7.800 55.100 8.200 55.200 ;
        RECT 15.000 55.100 15.400 55.200 ;
        RECT 33.400 55.100 33.800 55.200 ;
        RECT -2.600 54.800 33.800 55.100 ;
        RECT 34.200 53.100 34.600 53.200 ;
        RECT 35.000 53.100 35.400 53.200 ;
        RECT 34.200 52.800 35.400 53.100 ;
    END
  END B[0]
  PIN B[1]
    PORT
      LAYER metal1 ;
        RECT 8.800 46.900 9.200 47.000 ;
        RECT 8.700 46.600 9.200 46.900 ;
        RECT 18.100 46.800 18.600 47.200 ;
        RECT 5.400 45.800 5.800 46.600 ;
        RECT 8.700 46.200 9.000 46.600 ;
        RECT 18.000 46.400 18.400 46.800 ;
        RECT 8.600 45.800 9.000 46.200 ;
        RECT 11.000 45.400 11.400 46.200 ;
        RECT 26.200 44.400 26.600 45.200 ;
        RECT 10.200 34.400 10.600 35.200 ;
        RECT 16.000 34.200 16.400 34.600 ;
        RECT 12.600 33.800 13.000 34.200 ;
        RECT 14.200 34.100 14.600 34.200 ;
        RECT 15.800 34.100 16.300 34.200 ;
        RECT 14.200 33.800 16.300 34.100 ;
        RECT 12.600 33.200 12.900 33.800 ;
        RECT 12.600 32.400 13.000 33.200 ;
      LAYER via1 ;
        RECT 18.200 46.800 18.600 47.200 ;
        RECT 11.000 45.800 11.400 46.200 ;
        RECT 26.200 44.800 26.600 45.200 ;
        RECT 10.200 34.800 10.600 35.200 ;
      LAYER metal2 ;
        RECT 18.200 46.800 18.600 47.200 ;
        RECT 5.400 45.800 5.800 46.200 ;
        RECT 8.600 45.800 9.000 46.200 ;
        RECT 11.000 45.800 11.400 46.200 ;
        RECT 5.400 45.200 5.700 45.800 ;
        RECT 8.600 45.200 8.900 45.800 ;
        RECT 11.000 45.200 11.300 45.800 ;
        RECT 18.200 45.200 18.500 46.800 ;
        RECT 5.400 44.800 5.800 45.200 ;
        RECT 8.600 44.800 9.000 45.200 ;
        RECT 11.000 44.800 11.400 45.200 ;
        RECT 18.200 44.800 18.600 45.200 ;
        RECT 26.200 44.800 26.600 45.200 ;
        RECT 10.200 34.800 10.600 35.200 ;
        RECT 10.200 33.200 10.500 34.800 ;
        RECT 11.000 33.200 11.300 44.800 ;
        RECT 18.200 42.200 18.500 44.800 ;
        RECT 26.200 42.200 26.500 44.800 ;
        RECT 18.200 41.800 18.600 42.200 ;
        RECT 26.200 41.800 26.600 42.200 ;
        RECT 12.600 33.800 13.000 34.200 ;
        RECT 14.200 33.800 14.600 34.200 ;
        RECT 12.600 33.200 12.900 33.800 ;
        RECT 14.200 33.200 14.500 33.800 ;
        RECT 10.200 32.800 10.600 33.200 ;
        RECT 11.000 32.800 11.400 33.200 ;
        RECT 12.600 32.800 13.000 33.200 ;
        RECT 14.200 32.800 14.600 33.200 ;
      LAYER metal3 ;
        RECT -2.600 45.100 -2.200 45.200 ;
        RECT 5.400 45.100 5.800 45.200 ;
        RECT 8.600 45.100 9.000 45.200 ;
        RECT 11.000 45.100 11.400 45.200 ;
        RECT 18.200 45.100 18.600 45.200 ;
        RECT -2.600 44.800 18.600 45.100 ;
        RECT 18.200 42.100 18.600 42.200 ;
        RECT 26.200 42.100 26.600 42.200 ;
        RECT 18.200 41.800 26.600 42.100 ;
        RECT 10.200 33.100 10.600 33.200 ;
        RECT 11.000 33.100 11.400 33.200 ;
        RECT 12.600 33.100 13.000 33.200 ;
        RECT 14.200 33.100 14.600 33.200 ;
        RECT 10.200 32.800 14.600 33.100 ;
    END
  END B[1]
  PIN B[2]
    PORT
      LAYER metal1 ;
        RECT 26.200 32.400 26.600 33.200 ;
        RECT 25.400 26.800 25.900 27.200 ;
        RECT 25.600 26.400 26.000 26.800 ;
        RECT 6.200 14.100 6.600 14.200 ;
        RECT 7.000 14.100 7.400 14.200 ;
        RECT 6.200 13.800 7.800 14.100 ;
        RECT 7.400 13.600 7.800 13.800 ;
        RECT 24.600 13.400 25.000 14.200 ;
        RECT 9.400 7.800 9.800 8.600 ;
        RECT 23.000 7.800 23.400 8.600 ;
        RECT 5.000 7.100 5.800 7.200 ;
        RECT 6.200 7.100 6.600 7.200 ;
        RECT 4.700 7.000 6.600 7.100 ;
        RECT 3.600 6.800 6.600 7.000 ;
        RECT 3.600 6.700 5.000 6.800 ;
        RECT 3.600 6.600 4.000 6.700 ;
        RECT 6.200 6.400 6.600 6.800 ;
      LAYER via1 ;
        RECT 26.200 32.800 26.600 33.200 ;
        RECT 24.600 13.800 25.000 14.200 ;
        RECT 6.200 6.800 6.600 7.200 ;
      LAYER metal2 ;
        RECT 26.200 33.100 26.600 33.200 ;
        RECT 25.400 32.800 26.600 33.100 ;
        RECT 25.400 27.200 25.700 32.800 ;
        RECT 25.400 26.800 25.800 27.200 ;
        RECT 25.400 14.200 25.700 26.800 ;
        RECT 6.200 13.800 6.600 14.200 ;
        RECT 23.000 13.800 23.400 14.200 ;
        RECT 24.600 14.100 25.000 14.200 ;
        RECT 25.400 14.100 25.800 14.200 ;
        RECT 24.600 13.800 25.800 14.100 ;
        RECT 6.200 7.200 6.500 13.800 ;
        RECT 23.000 8.200 23.300 13.800 ;
        RECT 9.400 7.800 9.800 8.200 ;
        RECT 23.000 7.800 23.400 8.200 ;
        RECT 9.400 7.200 9.700 7.800 ;
        RECT 6.200 6.800 6.600 7.200 ;
        RECT 9.400 6.800 9.800 7.200 ;
      LAYER via2 ;
        RECT 25.400 13.800 25.800 14.200 ;
      LAYER metal3 ;
        RECT 6.200 14.100 6.600 14.200 ;
        RECT 23.000 14.100 23.400 14.200 ;
        RECT 25.400 14.100 25.800 14.200 ;
        RECT 6.200 13.800 25.800 14.100 ;
        RECT -2.600 7.100 -2.200 7.200 ;
        RECT 6.200 7.100 6.600 7.200 ;
        RECT 9.400 7.100 9.800 7.200 ;
        RECT -2.600 6.800 9.800 7.100 ;
    END
  END B[2]
  PIN B[3]
    PORT
      LAYER metal1 ;
        RECT 39.800 27.800 40.200 28.600 ;
        RECT 31.000 7.800 31.400 8.600 ;
        RECT 39.800 7.800 40.200 8.600 ;
        RECT 36.600 6.800 37.000 7.600 ;
        RECT 47.000 7.100 47.400 7.200 ;
        RECT 47.800 7.100 48.600 7.200 ;
        RECT 47.000 7.000 48.900 7.100 ;
        RECT 47.000 6.800 50.000 7.000 ;
        RECT 36.600 6.200 36.900 6.800 ;
        RECT 47.000 6.400 47.400 6.800 ;
        RECT 48.600 6.700 50.000 6.800 ;
        RECT 49.600 6.600 50.000 6.700 ;
        RECT 36.600 5.800 37.000 6.200 ;
      LAYER metal2 ;
        RECT 39.800 27.800 40.200 28.200 ;
        RECT 39.800 17.200 40.100 27.800 ;
        RECT 39.800 16.800 40.200 17.200 ;
        RECT 31.000 7.800 31.400 8.200 ;
        RECT 39.800 7.800 40.200 8.200 ;
        RECT 31.000 7.200 31.300 7.800 ;
        RECT 39.800 7.200 40.100 7.800 ;
        RECT 31.000 6.800 31.400 7.200 ;
        RECT 36.600 6.800 37.000 7.200 ;
        RECT 39.800 6.800 40.200 7.200 ;
        RECT 47.000 6.800 47.400 7.200 ;
        RECT 36.600 6.200 36.900 6.800 ;
        RECT 47.000 6.200 47.300 6.800 ;
        RECT 36.600 5.800 37.000 6.200 ;
        RECT 47.000 5.800 47.400 6.200 ;
        RECT 47.000 -1.800 47.300 5.800 ;
        RECT 47.000 -2.200 47.400 -1.800 ;
      LAYER metal3 ;
        RECT 39.800 16.800 40.200 17.200 ;
        RECT 39.800 16.200 40.100 16.800 ;
        RECT 39.800 15.800 40.200 16.200 ;
        RECT 31.000 7.100 31.400 7.200 ;
        RECT 36.600 7.100 37.000 7.200 ;
        RECT 39.800 7.100 40.200 7.200 ;
        RECT 31.000 6.800 40.200 7.100 ;
        RECT 39.800 6.100 40.100 6.800 ;
        RECT 47.000 6.100 47.400 6.200 ;
        RECT 39.800 5.800 47.400 6.100 ;
      LAYER via3 ;
        RECT 39.800 6.800 40.200 7.200 ;
      LAYER metal4 ;
        RECT 39.800 15.800 40.200 16.200 ;
        RECT 39.800 7.200 40.100 15.800 ;
        RECT 39.800 6.800 40.200 7.200 ;
    END
  END B[3]
  PIN B[4]
    PORT
      LAYER metal1 ;
        RECT 62.600 7.100 63.400 7.200 ;
        RECT 62.300 7.000 63.400 7.100 ;
        RECT 61.200 6.800 63.400 7.000 ;
        RECT 71.800 6.800 72.200 7.600 ;
        RECT 73.400 6.800 73.800 7.600 ;
        RECT 61.200 6.700 62.600 6.800 ;
        RECT 61.200 6.600 61.600 6.700 ;
        RECT 73.400 6.200 73.700 6.800 ;
        RECT 73.400 5.800 73.800 6.200 ;
      LAYER via1 ;
        RECT 63.000 6.800 63.400 7.200 ;
      LAYER metal2 ;
        RECT 63.000 6.800 63.400 7.200 ;
        RECT 71.800 7.100 72.200 7.200 ;
        RECT 72.600 7.100 73.000 7.200 ;
        RECT 71.800 6.800 73.000 7.100 ;
        RECT 73.400 6.800 73.800 7.200 ;
        RECT 63.000 5.200 63.300 6.800 ;
        RECT 71.800 5.200 72.100 6.800 ;
        RECT 73.400 6.200 73.700 6.800 ;
        RECT 73.400 5.800 73.800 6.200 ;
        RECT 63.000 4.800 63.400 5.200 ;
        RECT 71.800 4.800 72.200 5.200 ;
        RECT 63.000 -1.800 63.300 4.800 ;
        RECT 63.000 -2.200 63.400 -1.800 ;
      LAYER via2 ;
        RECT 72.600 6.800 73.000 7.200 ;
      LAYER metal3 ;
        RECT 72.600 7.100 73.000 7.200 ;
        RECT 73.400 7.100 73.800 7.200 ;
        RECT 72.600 6.800 73.800 7.100 ;
        RECT 63.000 5.100 63.400 5.200 ;
        RECT 71.800 5.100 72.200 5.200 ;
        RECT 63.000 4.800 72.200 5.100 ;
    END
  END B[4]
  PIN B[5]
    PORT
      LAYER metal1 ;
        RECT 72.600 34.100 73.000 34.200 ;
        RECT 72.200 33.800 73.000 34.100 ;
        RECT 72.200 33.600 72.600 33.800 ;
        RECT 75.000 33.400 75.400 34.200 ;
        RECT 91.800 32.400 92.200 33.200 ;
        RECT 95.400 7.100 96.200 7.200 ;
        RECT 97.400 7.100 97.800 7.200 ;
        RECT 95.100 7.000 97.800 7.100 ;
        RECT 94.000 6.800 97.800 7.000 ;
        RECT 94.000 6.700 95.400 6.800 ;
        RECT 94.000 6.600 94.400 6.700 ;
      LAYER via1 ;
        RECT 72.600 33.800 73.000 34.200 ;
        RECT 75.000 33.800 75.400 34.200 ;
        RECT 91.800 32.800 92.200 33.200 ;
        RECT 97.400 6.800 97.800 7.200 ;
      LAYER metal2 ;
        RECT 72.600 33.800 73.000 34.200 ;
        RECT 75.000 33.800 75.400 34.200 ;
        RECT 72.600 33.200 72.900 33.800 ;
        RECT 75.000 33.200 75.300 33.800 ;
        RECT 72.600 32.800 73.000 33.200 ;
        RECT 75.000 32.800 75.400 33.200 ;
        RECT 91.800 33.100 92.200 33.200 ;
        RECT 92.600 33.100 93.000 33.200 ;
        RECT 91.800 32.800 93.000 33.100 ;
        RECT 97.400 25.800 97.800 26.200 ;
        RECT 97.400 7.200 97.700 25.800 ;
        RECT 97.400 6.800 97.800 7.200 ;
      LAYER via2 ;
        RECT 92.600 32.800 93.000 33.200 ;
      LAYER metal3 ;
        RECT 72.600 33.100 73.000 33.200 ;
        RECT 75.000 33.100 75.400 33.200 ;
        RECT 75.800 33.100 76.200 33.200 ;
        RECT 72.600 32.800 76.200 33.100 ;
        RECT 91.800 33.100 92.200 33.200 ;
        RECT 92.600 33.100 93.000 33.200 ;
        RECT 91.800 32.800 93.000 33.100 ;
        RECT 97.400 26.100 97.800 26.200 ;
        RECT 100.600 26.100 101.000 26.200 ;
        RECT 97.400 25.800 101.000 26.100 ;
      LAYER via3 ;
        RECT 75.800 32.800 76.200 33.200 ;
      LAYER metal4 ;
        RECT 75.000 33.100 75.400 33.200 ;
        RECT 75.800 33.100 76.200 33.200 ;
        RECT 75.000 32.800 76.200 33.100 ;
        RECT 91.800 33.100 92.200 33.200 ;
        RECT 92.600 33.100 93.000 33.200 ;
        RECT 91.800 32.800 93.000 33.100 ;
        RECT 97.400 32.800 97.800 33.200 ;
        RECT 97.400 26.200 97.700 32.800 ;
        RECT 97.400 25.800 97.800 26.200 ;
      LAYER via4 ;
        RECT 92.600 32.800 93.000 33.200 ;
      LAYER metal5 ;
        RECT 75.000 33.100 75.400 33.200 ;
        RECT 92.600 33.100 93.000 33.200 ;
        RECT 97.400 33.100 97.800 33.200 ;
        RECT 75.000 32.800 97.800 33.100 ;
    END
  END B[5]
  PIN B[6]
    PORT
      LAYER metal1 ;
        RECT 78.200 67.800 78.600 68.600 ;
        RECT 78.200 52.400 78.600 53.200 ;
        RECT 90.200 52.400 90.600 53.200 ;
      LAYER via1 ;
        RECT 78.200 52.800 78.600 53.200 ;
        RECT 90.200 52.800 90.600 53.200 ;
      LAYER metal2 ;
        RECT 78.200 68.100 78.600 68.200 ;
        RECT 79.000 68.100 79.400 68.200 ;
        RECT 78.200 67.800 79.400 68.100 ;
        RECT 78.200 53.800 78.600 54.200 ;
        RECT 90.200 53.800 90.600 54.200 ;
        RECT 78.200 53.200 78.500 53.800 ;
        RECT 90.200 53.200 90.500 53.800 ;
        RECT 78.200 52.800 78.600 53.200 ;
        RECT 90.200 52.800 90.600 53.200 ;
      LAYER via2 ;
        RECT 79.000 67.800 79.400 68.200 ;
      LAYER metal3 ;
        RECT 78.200 68.100 78.600 68.200 ;
        RECT 79.000 68.100 79.400 68.200 ;
        RECT 78.200 67.800 79.400 68.100 ;
        RECT 97.400 56.100 97.800 56.200 ;
        RECT 100.600 56.100 101.000 56.200 ;
        RECT 97.400 55.800 101.000 56.100 ;
        RECT 78.200 54.100 78.600 54.200 ;
        RECT 90.200 54.100 90.600 54.200 ;
        RECT 97.400 54.100 97.800 54.200 ;
        RECT 78.200 53.800 97.800 54.100 ;
        RECT 78.200 53.200 78.500 53.800 ;
        RECT 78.200 52.800 78.600 53.200 ;
      LAYER via3 ;
        RECT 97.400 53.800 97.800 54.200 ;
      LAYER metal4 ;
        RECT 78.200 67.800 78.600 68.200 ;
        RECT 78.200 53.200 78.500 67.800 ;
        RECT 97.400 55.800 97.800 56.200 ;
        RECT 97.400 54.200 97.700 55.800 ;
        RECT 97.400 53.800 97.800 54.200 ;
        RECT 78.200 52.800 78.600 53.200 ;
    END
  END B[6]
  PIN B[7]
    PORT
      LAYER metal1 ;
        RECT 43.800 73.800 44.200 74.200 ;
        RECT 43.800 73.200 44.100 73.800 ;
        RECT 43.800 72.400 44.200 73.200 ;
        RECT 48.600 72.400 49.000 73.200 ;
      LAYER via1 ;
        RECT 48.600 72.800 49.000 73.200 ;
      LAYER metal2 ;
        RECT 47.000 82.800 47.400 83.200 ;
        RECT 43.800 73.800 44.200 74.200 ;
        RECT 43.800 73.200 44.100 73.800 ;
        RECT 47.000 73.200 47.300 82.800 ;
        RECT 43.800 72.800 44.200 73.200 ;
        RECT 47.000 72.800 47.400 73.200 ;
        RECT 47.800 73.100 48.200 73.200 ;
        RECT 48.600 73.100 49.000 73.200 ;
        RECT 47.800 72.800 49.000 73.100 ;
      LAYER metal3 ;
        RECT 43.800 73.100 44.200 73.200 ;
        RECT 47.000 73.100 47.400 73.200 ;
        RECT 47.800 73.100 48.200 73.200 ;
        RECT 43.800 72.800 48.200 73.100 ;
    END
  END B[7]
  PIN opcode[0]
    PORT
      LAYER metal1 ;
        RECT 8.600 73.400 9.000 74.200 ;
        RECT 15.000 74.100 15.400 74.200 ;
        RECT 14.200 73.800 15.400 74.100 ;
        RECT 14.200 73.200 14.500 73.800 ;
        RECT 15.000 73.400 15.400 73.800 ;
        RECT 4.600 72.400 5.000 73.200 ;
        RECT 14.200 72.400 14.600 73.200 ;
        RECT 17.400 72.400 17.800 73.200 ;
      LAYER via1 ;
        RECT 8.600 73.800 9.000 74.200 ;
        RECT 15.000 73.800 15.400 74.200 ;
        RECT 4.600 72.800 5.000 73.200 ;
        RECT 17.400 72.800 17.800 73.200 ;
      LAYER metal2 ;
        RECT 4.600 73.800 5.000 74.200 ;
        RECT 8.600 74.100 9.000 74.200 ;
        RECT 9.400 74.100 9.800 74.200 ;
        RECT 8.600 73.800 9.800 74.100 ;
        RECT 15.000 74.100 15.400 74.200 ;
        RECT 15.800 74.100 16.200 74.200 ;
        RECT 15.000 73.800 16.200 74.100 ;
        RECT 17.400 73.800 17.800 74.200 ;
        RECT 4.600 73.200 4.900 73.800 ;
        RECT 17.400 73.200 17.700 73.800 ;
        RECT 4.600 72.800 5.000 73.200 ;
        RECT 17.400 72.800 17.800 73.200 ;
      LAYER via2 ;
        RECT 9.400 73.800 9.800 74.200 ;
        RECT 15.800 73.800 16.200 74.200 ;
      LAYER metal3 ;
        RECT -2.600 74.100 -2.200 74.200 ;
        RECT 4.600 74.100 5.000 74.200 ;
        RECT 9.400 74.100 9.800 74.200 ;
        RECT 15.800 74.100 16.200 74.200 ;
        RECT 17.400 74.100 17.800 74.200 ;
        RECT -2.600 73.800 17.800 74.100 ;
    END
  END opcode[0]
  PIN opcode[1]
    PORT
      LAYER metal1 ;
        RECT 10.200 76.100 10.600 77.200 ;
        RECT 11.000 76.100 11.400 76.200 ;
        RECT 10.200 75.800 11.400 76.100 ;
        RECT 12.600 74.800 13.000 75.600 ;
        RECT 7.800 73.400 8.200 74.200 ;
        RECT 11.000 72.400 11.400 73.200 ;
      LAYER via1 ;
        RECT 10.200 76.800 10.600 77.200 ;
        RECT 11.000 75.800 11.400 76.200 ;
        RECT 7.800 73.800 8.200 74.200 ;
        RECT 11.000 72.800 11.400 73.200 ;
      LAYER metal2 ;
        RECT 10.200 82.800 10.600 83.200 ;
        RECT 10.200 77.200 10.500 82.800 ;
        RECT 10.200 76.800 10.600 77.200 ;
        RECT 11.000 75.800 11.400 76.200 ;
        RECT 7.800 73.800 8.200 74.200 ;
        RECT 7.800 73.200 8.100 73.800 ;
        RECT 11.000 73.200 11.300 75.800 ;
        RECT 12.600 74.800 13.000 75.200 ;
        RECT 12.600 73.200 12.900 74.800 ;
        RECT 7.800 72.800 8.200 73.200 ;
        RECT 11.000 73.100 11.400 73.200 ;
        RECT 11.800 73.100 12.200 73.200 ;
        RECT 11.000 72.800 12.200 73.100 ;
        RECT 12.600 72.800 13.000 73.200 ;
      LAYER via2 ;
        RECT 11.800 72.800 12.200 73.200 ;
      LAYER metal3 ;
        RECT 7.800 73.100 8.200 73.200 ;
        RECT 11.800 73.100 12.200 73.200 ;
        RECT 12.600 73.100 13.000 73.200 ;
        RECT 7.800 72.800 13.000 73.100 ;
    END
  END opcode[1]
  PIN opcode[2]
    PORT
      LAYER metal1 ;
        RECT 23.800 74.800 24.200 75.200 ;
        RECT 32.600 74.800 33.000 75.600 ;
        RECT 23.800 74.400 24.100 74.800 ;
        RECT 23.600 74.100 24.100 74.400 ;
        RECT 23.600 74.000 24.000 74.100 ;
        RECT 25.400 73.400 25.800 74.200 ;
        RECT 39.800 72.800 40.200 73.200 ;
        RECT 39.900 72.400 40.300 72.800 ;
      LAYER via1 ;
        RECT 25.400 73.800 25.800 74.200 ;
      LAYER metal2 ;
        RECT 32.600 82.800 33.000 83.200 ;
        RECT 32.600 75.200 32.900 82.800 ;
        RECT 23.800 74.800 24.200 75.200 ;
        RECT 32.600 74.800 33.000 75.200 ;
        RECT 23.800 74.200 24.100 74.800 ;
        RECT 32.600 74.200 32.900 74.800 ;
        RECT 23.800 73.800 24.200 74.200 ;
        RECT 24.600 74.100 25.000 74.200 ;
        RECT 25.400 74.100 25.800 74.200 ;
        RECT 24.600 73.800 25.800 74.100 ;
        RECT 32.600 73.800 33.000 74.200 ;
        RECT 39.800 73.800 40.200 74.200 ;
        RECT 39.800 73.200 40.100 73.800 ;
        RECT 39.800 72.800 40.200 73.200 ;
      LAYER metal3 ;
        RECT 23.800 74.100 24.200 74.200 ;
        RECT 24.600 74.100 25.000 74.200 ;
        RECT 32.600 74.100 33.000 74.200 ;
        RECT 39.800 74.100 40.200 74.200 ;
        RECT 23.800 73.800 40.200 74.100 ;
    END
  END opcode[2]
  PIN opcode[3]
    PORT
      LAYER metal1 ;
        RECT 35.800 75.100 36.200 75.200 ;
        RECT 36.600 75.100 37.000 76.200 ;
        RECT 35.800 74.800 37.000 75.100 ;
        RECT 30.200 72.400 30.600 73.200 ;
        RECT 34.200 72.400 34.600 73.200 ;
        RECT 40.600 67.800 41.000 68.600 ;
      LAYER via1 ;
        RECT 30.200 72.800 30.600 73.200 ;
        RECT 34.200 72.800 34.600 73.200 ;
      LAYER metal2 ;
        RECT 35.000 83.100 35.400 83.200 ;
        RECT 35.000 82.800 36.100 83.100 ;
        RECT 35.800 75.200 36.100 82.800 ;
        RECT 30.200 74.800 30.600 75.200 ;
        RECT 34.200 74.800 34.600 75.200 ;
        RECT 35.800 74.800 36.200 75.200 ;
        RECT 40.600 74.800 41.000 75.200 ;
        RECT 30.200 73.200 30.500 74.800 ;
        RECT 34.200 73.200 34.500 74.800 ;
        RECT 30.200 72.800 30.600 73.200 ;
        RECT 34.200 72.800 34.600 73.200 ;
        RECT 40.600 68.200 40.900 74.800 ;
        RECT 40.600 67.800 41.000 68.200 ;
      LAYER metal3 ;
        RECT 30.200 75.100 30.600 75.200 ;
        RECT 34.200 75.100 34.600 75.200 ;
        RECT 35.800 75.100 36.200 75.200 ;
        RECT 40.600 75.100 41.000 75.200 ;
        RECT 30.200 74.800 41.000 75.100 ;
    END
  END opcode[3]
  PIN result[0]
    PORT
      LAYER metal1 ;
        RECT 57.400 6.200 57.800 9.900 ;
        RECT 57.500 5.100 57.800 6.200 ;
        RECT 57.400 1.100 57.800 5.100 ;
      LAYER via1 ;
        RECT 57.400 1.800 57.800 2.200 ;
      LAYER metal2 ;
        RECT 57.400 1.800 57.800 2.200 ;
        RECT 56.600 -1.900 57.000 -1.800 ;
        RECT 57.400 -1.900 57.700 1.800 ;
        RECT 56.600 -2.200 57.700 -1.900 ;
    END
  END result[0]
  PIN result[1]
    PORT
      LAYER metal1 ;
        RECT 0.600 75.900 1.000 79.900 ;
        RECT 0.600 74.800 0.900 75.900 ;
        RECT 0.600 71.100 1.000 74.800 ;
      LAYER via1 ;
        RECT 0.600 76.800 1.000 77.200 ;
      LAYER metal2 ;
        RECT 0.600 76.800 1.000 77.200 ;
        RECT 0.600 76.200 0.900 76.800 ;
        RECT 0.600 75.800 1.000 76.200 ;
      LAYER metal3 ;
        RECT -2.600 76.100 -2.200 76.200 ;
        RECT 0.600 76.100 1.000 76.200 ;
        RECT -2.600 75.800 1.000 76.100 ;
    END
  END result[1]
  PIN result[2]
    PORT
      LAYER metal1 ;
        RECT 0.600 26.200 1.000 29.900 ;
        RECT 0.600 25.100 0.900 26.200 ;
        RECT 0.600 21.100 1.000 25.100 ;
      LAYER via1 ;
        RECT 0.600 23.800 1.000 24.200 ;
      LAYER metal2 ;
        RECT 0.600 24.800 1.000 25.200 ;
        RECT 0.600 24.200 0.900 24.800 ;
        RECT 0.600 23.800 1.000 24.200 ;
      LAYER metal3 ;
        RECT -2.600 25.100 -2.200 25.200 ;
        RECT 0.600 25.100 1.000 25.200 ;
        RECT -2.600 24.800 1.000 25.100 ;
    END
  END result[2]
  PIN result[3]
    PORT
      LAYER metal1 ;
        RECT 55.000 6.200 55.400 9.900 ;
        RECT 55.100 5.100 55.400 6.200 ;
        RECT 55.000 1.100 55.400 5.100 ;
      LAYER via1 ;
        RECT 55.000 1.800 55.400 2.200 ;
      LAYER metal2 ;
        RECT 55.000 1.800 55.400 2.200 ;
        RECT 54.200 -1.900 54.600 -1.800 ;
        RECT 55.000 -1.900 55.300 1.800 ;
        RECT 54.200 -2.200 55.300 -1.900 ;
    END
  END result[3]
  PIN result[4]
    PORT
      LAYER metal1 ;
        RECT 94.200 75.900 94.600 79.900 ;
        RECT 94.300 74.800 94.600 75.900 ;
        RECT 94.200 71.100 94.600 74.800 ;
      LAYER via1 ;
        RECT 94.200 71.800 94.600 72.200 ;
      LAYER metal2 ;
        RECT 94.200 71.800 94.600 72.200 ;
        RECT 94.200 68.200 94.500 71.800 ;
        RECT 94.200 67.800 94.600 68.200 ;
        RECT 93.400 0.800 93.800 1.200 ;
        RECT 93.400 -1.800 93.700 0.800 ;
        RECT 93.400 -2.200 93.800 -1.800 ;
      LAYER metal3 ;
        RECT 93.400 68.100 93.800 68.200 ;
        RECT 94.200 68.100 94.600 68.200 ;
        RECT 93.400 67.800 94.600 68.100 ;
        RECT 93.400 1.100 93.800 1.200 ;
        RECT 94.200 1.100 94.600 1.200 ;
        RECT 93.400 0.800 94.600 1.100 ;
      LAYER via3 ;
        RECT 94.200 0.800 94.600 1.200 ;
      LAYER metal4 ;
        RECT 93.400 67.800 93.800 68.200 ;
        RECT 93.400 1.100 93.700 67.800 ;
        RECT 94.200 1.100 94.600 1.200 ;
        RECT 93.400 0.800 94.600 1.100 ;
    END
  END result[4]
  PIN result[5]
    PORT
      LAYER metal1 ;
        RECT 87.000 6.200 87.400 9.900 ;
        RECT 87.000 5.100 87.300 6.200 ;
        RECT 87.000 1.100 87.400 5.100 ;
      LAYER via1 ;
        RECT 87.000 1.800 87.400 2.200 ;
      LAYER metal2 ;
        RECT 87.000 1.800 87.400 2.200 ;
        RECT 87.000 -1.900 87.300 1.800 ;
        RECT 87.800 -1.900 88.200 -1.800 ;
        RECT 87.000 -2.200 88.200 -1.900 ;
    END
  END result[5]
  PIN result[6]
    PORT
      LAYER metal1 ;
        RECT 94.200 46.200 94.600 49.900 ;
        RECT 94.300 45.100 94.600 46.200 ;
        RECT 94.200 41.100 94.600 45.100 ;
      LAYER via1 ;
        RECT 94.200 43.800 94.600 44.200 ;
      LAYER metal2 ;
        RECT 94.200 44.800 94.600 45.200 ;
        RECT 94.200 44.200 94.500 44.800 ;
        RECT 94.200 43.800 94.600 44.200 ;
      LAYER metal3 ;
        RECT 94.200 45.100 94.600 45.200 ;
        RECT 100.600 45.100 101.000 45.200 ;
        RECT 94.200 44.800 101.000 45.100 ;
    END
  END result[6]
  PIN result[7]
    PORT
      LAYER metal1 ;
        RECT 95.000 75.900 95.400 79.900 ;
        RECT 95.000 74.800 95.300 75.900 ;
        RECT 95.000 71.100 95.400 74.800 ;
      LAYER via1 ;
        RECT 95.000 78.800 95.400 79.200 ;
      LAYER metal2 ;
        RECT 95.800 83.100 96.200 83.200 ;
        RECT 95.000 82.800 96.200 83.100 ;
        RECT 95.000 79.200 95.300 82.800 ;
        RECT 95.000 78.800 95.400 79.200 ;
    END
  END result[7]
  PIN overflow
    PORT
      LAYER metal1 ;
        RECT 89.400 75.900 89.800 79.900 ;
        RECT 89.500 74.800 89.800 75.900 ;
        RECT 89.400 71.100 89.800 74.800 ;
      LAYER via1 ;
        RECT 89.400 78.800 89.800 79.200 ;
      LAYER metal2 ;
        RECT 88.600 83.100 89.000 83.200 ;
        RECT 88.600 82.800 89.700 83.100 ;
        RECT 89.400 79.200 89.700 82.800 ;
        RECT 89.400 78.800 89.800 79.200 ;
    END
  END overflow
  PIN negative
    PORT
      LAYER metal1 ;
        RECT 91.800 75.900 92.200 79.900 ;
        RECT 91.900 74.800 92.200 75.900 ;
        RECT 91.800 71.100 92.200 74.800 ;
      LAYER via1 ;
        RECT 91.800 78.800 92.200 79.200 ;
      LAYER metal2 ;
        RECT 91.000 83.100 91.400 83.200 ;
        RECT 91.000 82.800 92.100 83.100 ;
        RECT 91.800 79.200 92.100 82.800 ;
        RECT 91.800 78.800 92.200 79.200 ;
    END
  END negative
  PIN zero
    PORT
      LAYER metal1 ;
        RECT 94.200 55.900 94.600 59.900 ;
        RECT 94.300 54.800 94.600 55.900 ;
        RECT 94.200 51.100 94.600 54.800 ;
      LAYER via1 ;
        RECT 94.200 58.800 94.600 59.200 ;
      LAYER metal2 ;
        RECT 94.200 59.800 94.600 60.200 ;
        RECT 94.200 59.200 94.500 59.800 ;
        RECT 94.200 58.800 94.600 59.200 ;
      LAYER metal3 ;
        RECT 94.200 60.100 94.600 60.200 ;
        RECT 100.600 60.100 101.000 60.200 ;
        RECT 94.200 59.800 101.000 60.100 ;
    END
  END zero
  OBS
      LAYER metal1 ;
        RECT 2.200 76.200 2.600 79.900 ;
        RECT 1.500 75.900 2.600 76.200 ;
        RECT 1.500 75.600 1.800 75.900 ;
        RECT 1.200 75.200 1.800 75.600 ;
        RECT 1.500 73.700 1.800 75.200 ;
        RECT 2.200 75.100 2.600 75.200 ;
        RECT 3.000 75.100 3.400 79.900 ;
        RECT 2.200 74.800 3.400 75.100 ;
        RECT 2.200 74.400 2.600 74.800 ;
        RECT 1.500 73.400 2.600 73.700 ;
        RECT 2.200 71.100 2.600 73.400 ;
        RECT 3.000 71.100 3.400 74.800 ;
        RECT 5.400 76.100 5.800 79.900 ;
        RECT 6.200 76.100 6.600 76.600 ;
        RECT 5.400 75.800 6.600 76.100 ;
        RECT 3.800 72.400 4.200 73.200 ;
        RECT 5.400 71.100 5.800 75.800 ;
        RECT 7.000 73.100 7.400 79.900 ;
        RECT 6.500 72.800 7.400 73.100 ;
        RECT 9.400 73.100 9.800 79.900 ;
        RECT 9.400 72.800 10.300 73.100 ;
        RECT 6.500 72.200 6.900 72.800 ;
        RECT 9.900 72.200 10.300 72.800 ;
        RECT 6.500 71.800 7.400 72.200 ;
        RECT 9.900 71.800 10.600 72.200 ;
        RECT 6.500 71.100 6.900 71.800 ;
        RECT 9.900 71.100 10.300 71.800 ;
        RECT 11.800 71.100 12.200 79.900 ;
        RECT 12.900 77.200 13.300 79.900 ;
        RECT 12.900 76.800 13.800 77.200 ;
        RECT 12.900 76.300 13.300 76.800 ;
        RECT 12.900 75.900 13.800 76.300 ;
        RECT 13.400 74.200 13.700 75.900 ;
        RECT 13.400 73.800 13.800 74.200 ;
        RECT 13.400 72.100 13.700 73.800 ;
        RECT 15.800 73.100 16.200 79.900 ;
        RECT 16.600 75.800 17.000 76.600 ;
        RECT 18.700 76.300 19.100 79.900 ;
        RECT 18.200 75.900 19.100 76.300 ;
        RECT 18.300 74.200 18.600 75.900 ;
        RECT 19.000 74.800 19.400 75.600 ;
        RECT 18.200 74.100 18.600 74.200 ;
        RECT 19.800 74.100 20.200 74.200 ;
        RECT 18.200 73.800 20.200 74.100 ;
        RECT 15.800 72.800 16.700 73.100 ;
        RECT 16.300 72.200 16.700 72.800 ;
        RECT 13.400 71.100 13.800 72.100 ;
        RECT 16.300 71.800 17.000 72.200 ;
        RECT 18.300 72.100 18.600 73.800 ;
        RECT 19.800 73.400 20.200 73.800 ;
        RECT 20.600 73.100 21.000 79.900 ;
        RECT 21.400 76.100 21.800 76.600 ;
        RECT 22.200 76.100 22.600 79.900 ;
        RECT 21.400 75.900 22.600 76.100 ;
        RECT 23.800 77.900 24.200 79.900 ;
        RECT 21.400 75.800 22.500 75.900 ;
        RECT 23.800 75.800 24.100 77.900 ;
        RECT 22.200 75.200 22.500 75.800 ;
        RECT 22.900 75.500 24.100 75.800 ;
        RECT 22.200 74.800 22.600 75.200 ;
        RECT 22.200 73.100 22.500 74.800 ;
        RECT 22.900 73.800 23.200 75.500 ;
        RECT 25.400 75.100 25.800 75.200 ;
        RECT 24.600 74.800 25.800 75.100 ;
        RECT 24.600 73.800 25.000 74.800 ;
        RECT 22.800 73.700 23.200 73.800 ;
        RECT 22.800 73.500 24.300 73.700 ;
        RECT 22.800 73.400 24.900 73.500 ;
        RECT 24.000 73.200 24.900 73.400 ;
        RECT 24.600 73.100 24.900 73.200 ;
        RECT 26.200 73.100 26.600 79.900 ;
        RECT 27.000 76.100 27.400 76.600 ;
        RECT 29.400 76.100 29.800 79.900 ;
        RECT 27.000 75.800 29.800 76.100 ;
        RECT 20.600 72.800 21.500 73.100 ;
        RECT 16.300 71.100 16.700 71.800 ;
        RECT 18.200 71.100 18.600 72.100 ;
        RECT 21.100 72.200 21.500 72.800 ;
        RECT 22.200 72.600 22.900 73.100 ;
        RECT 21.100 71.800 21.800 72.200 ;
        RECT 21.100 71.100 21.500 71.800 ;
        RECT 22.500 71.100 22.900 72.600 ;
        RECT 24.600 71.100 25.000 73.100 ;
        RECT 26.200 72.800 27.100 73.100 ;
        RECT 26.700 72.200 27.100 72.800 ;
        RECT 26.200 71.800 27.100 72.200 ;
        RECT 26.700 71.100 27.100 71.800 ;
        RECT 29.400 71.100 29.800 75.800 ;
        RECT 31.000 71.100 31.400 79.900 ;
        RECT 32.900 76.300 33.300 79.900 ;
        RECT 32.900 75.900 33.800 76.300 ;
        RECT 33.400 74.200 33.700 75.900 ;
        RECT 31.800 74.100 32.200 74.200 ;
        RECT 33.400 74.100 33.800 74.200 ;
        RECT 31.800 73.800 33.800 74.100 ;
        RECT 31.800 73.400 32.200 73.800 ;
        RECT 33.400 72.100 33.700 73.800 ;
        RECT 33.400 71.100 33.800 72.100 ;
        RECT 35.000 71.100 35.400 79.900 ;
        RECT 37.400 77.900 37.800 79.900 ;
        RECT 37.500 77.800 37.800 77.900 ;
        RECT 39.000 77.900 39.400 79.900 ;
        RECT 39.000 77.800 39.300 77.900 ;
        RECT 37.500 77.500 39.300 77.800 ;
        RECT 38.200 76.400 38.600 77.200 ;
        RECT 39.000 76.200 39.300 77.500 ;
        RECT 39.000 75.800 39.400 76.200 ;
        RECT 39.800 75.900 40.200 79.900 ;
        RECT 40.600 76.200 41.000 79.900 ;
        RECT 42.200 76.200 42.600 79.900 ;
        RECT 40.600 75.900 42.600 76.200 ;
        RECT 37.400 74.800 38.200 75.200 ;
        RECT 39.000 74.200 39.300 75.800 ;
        RECT 39.900 75.200 40.200 75.900 ;
        RECT 39.800 74.900 41.000 75.200 ;
        RECT 39.800 74.800 40.200 74.900 ;
        RECT 35.800 73.400 36.200 74.200 ;
        RECT 38.500 74.100 39.300 74.200 ;
        RECT 38.400 73.900 39.300 74.100 ;
        RECT 38.400 72.200 38.800 73.900 ;
        RECT 40.700 73.100 41.000 74.900 ;
        RECT 43.000 75.100 43.400 79.900 ;
        RECT 45.900 76.300 46.300 79.900 ;
        RECT 45.400 75.900 46.300 76.300 ;
        RECT 44.600 75.100 45.000 75.200 ;
        RECT 43.000 74.800 45.000 75.100 ;
        RECT 41.400 74.100 41.800 74.600 ;
        RECT 43.000 74.100 43.400 74.800 ;
        RECT 45.500 74.200 45.800 75.900 ;
        RECT 46.200 75.100 46.600 75.600 ;
        RECT 47.000 75.100 47.400 79.900 ;
        RECT 49.900 76.300 50.300 79.900 ;
        RECT 49.400 75.900 50.300 76.300 ;
        RECT 51.300 76.300 51.700 79.900 ;
        RECT 51.300 75.900 52.200 76.300 ;
        RECT 46.200 74.800 47.400 75.100 ;
        RECT 41.400 73.800 43.400 74.100 ;
        RECT 45.400 73.800 45.800 74.200 ;
        RECT 38.400 71.800 39.400 72.200 ;
        RECT 38.400 71.100 38.800 71.800 ;
        RECT 40.600 71.100 41.000 73.100 ;
        RECT 43.000 71.100 43.400 73.800 ;
        RECT 44.600 72.400 45.000 73.200 ;
        RECT 45.500 72.200 45.800 73.800 ;
        RECT 45.400 71.100 45.800 72.200 ;
        RECT 47.000 71.100 47.400 74.800 ;
        RECT 49.500 74.200 49.800 75.900 ;
        RECT 51.000 74.800 51.400 75.600 ;
        RECT 49.400 73.800 49.800 74.200 ;
        RECT 49.500 73.200 49.800 73.800 ;
        RECT 49.400 72.800 49.800 73.200 ;
        RECT 49.500 72.100 49.800 72.800 ;
        RECT 49.400 71.100 49.800 72.100 ;
        RECT 51.800 74.200 52.100 75.900 ;
        RECT 51.800 74.100 52.200 74.200 ;
        RECT 53.400 74.100 53.800 74.200 ;
        RECT 51.800 73.800 53.800 74.100 ;
        RECT 51.800 72.100 52.100 73.800 ;
        RECT 53.400 73.400 53.800 73.800 ;
        RECT 54.200 74.100 54.600 79.900 ;
        RECT 55.900 79.600 57.700 79.900 ;
        RECT 55.900 79.500 56.200 79.600 ;
        RECT 55.800 76.500 56.200 79.500 ;
        RECT 57.400 79.500 57.700 79.600 ;
        RECT 58.200 79.600 60.200 79.900 ;
        RECT 56.600 76.500 57.000 79.300 ;
        RECT 57.400 76.700 57.800 79.500 ;
        RECT 58.200 77.000 58.600 79.600 ;
        RECT 59.000 76.900 59.400 79.300 ;
        RECT 59.800 76.900 60.200 79.600 ;
        RECT 59.000 76.700 59.300 76.900 ;
        RECT 57.400 76.500 59.300 76.700 ;
        RECT 56.700 76.200 57.000 76.500 ;
        RECT 57.500 76.400 59.300 76.500 ;
        RECT 59.900 76.600 60.200 76.900 ;
        RECT 61.400 76.900 61.800 79.900 ;
        RECT 61.400 76.600 61.700 76.900 ;
        RECT 59.900 76.300 61.700 76.600 ;
        RECT 56.600 76.100 57.000 76.200 ;
        RECT 56.600 75.800 58.300 76.100 ;
        RECT 62.200 75.900 62.600 79.900 ;
        RECT 63.000 76.200 63.400 79.900 ;
        RECT 64.600 76.200 65.000 79.900 ;
        RECT 65.800 76.800 66.200 77.200 ;
        RECT 65.800 76.200 66.100 76.800 ;
        RECT 66.500 76.200 66.900 79.900 ;
        RECT 71.000 77.800 71.400 79.900 ;
        RECT 72.600 77.900 73.000 79.900 ;
        RECT 72.600 77.800 72.900 77.900 ;
        RECT 71.100 77.500 72.900 77.800 ;
        RECT 71.800 76.400 72.200 77.200 ;
        RECT 72.600 76.200 72.900 77.500 ;
        RECT 63.000 75.900 65.000 76.200 ;
        RECT 65.400 75.900 66.100 76.200 ;
        RECT 66.400 75.900 66.900 76.200 ;
        RECT 55.000 74.100 55.400 74.200 ;
        RECT 54.200 73.800 55.400 74.100 ;
        RECT 52.600 72.400 53.000 73.200 ;
        RECT 51.800 71.100 52.200 72.100 ;
        RECT 54.200 71.100 54.600 73.800 ;
        RECT 58.000 72.500 58.300 75.800 ;
        RECT 62.300 75.200 62.600 75.900 ;
        RECT 65.400 75.800 65.800 75.900 ;
        RECT 64.200 75.200 64.600 75.400 ;
        RECT 58.600 75.100 59.400 75.200 ;
        RECT 61.400 75.100 61.800 75.200 ;
        RECT 58.600 74.800 61.800 75.100 ;
        RECT 62.200 74.900 63.400 75.200 ;
        RECT 64.200 74.900 65.000 75.200 ;
        RECT 62.200 74.800 62.600 74.900 ;
        RECT 63.100 74.100 63.400 74.900 ;
        RECT 64.600 74.800 65.000 74.900 ;
        RECT 60.600 73.800 63.400 74.100 ;
        RECT 63.800 74.100 64.200 74.600 ;
        RECT 66.400 74.200 66.700 75.900 ;
        RECT 70.200 75.400 70.600 76.200 ;
        RECT 72.600 75.800 73.000 76.200 ;
        RECT 67.000 74.400 67.400 75.200 ;
        RECT 71.000 74.800 71.800 75.200 ;
        RECT 72.600 74.200 72.900 75.800 ;
        RECT 65.400 74.100 66.700 74.200 ;
        RECT 67.800 74.100 68.200 74.200 ;
        RECT 72.100 74.100 72.900 74.200 ;
        RECT 63.800 73.800 66.700 74.100 ;
        RECT 67.400 73.800 68.200 74.100 ;
        RECT 72.000 73.900 72.900 74.100 ;
        RECT 73.400 75.100 73.800 79.900 ;
        RECT 75.000 77.900 75.400 79.900 ;
        RECT 75.100 77.800 75.400 77.900 ;
        RECT 76.600 77.900 77.000 79.900 ;
        RECT 76.600 77.800 76.900 77.900 ;
        RECT 75.100 77.500 76.900 77.800 ;
        RECT 75.100 76.200 75.400 77.500 ;
        RECT 75.800 76.400 76.200 77.200 ;
        RECT 78.200 76.200 78.600 79.900 ;
        RECT 79.800 76.200 80.200 79.900 ;
        RECT 75.000 75.800 75.400 76.200 ;
        RECT 74.200 75.100 74.600 75.200 ;
        RECT 73.400 74.800 74.600 75.100 ;
        RECT 60.600 73.200 60.900 73.800 ;
        RECT 60.100 72.800 61.000 73.200 ;
        RECT 62.200 72.800 62.600 73.200 ;
        RECT 63.100 73.100 63.400 73.800 ;
        RECT 65.500 73.100 65.800 73.800 ;
        RECT 67.400 73.600 67.800 73.800 ;
        RECT 66.300 73.100 68.100 73.300 ;
        RECT 58.000 72.200 60.000 72.500 ;
        RECT 62.300 72.400 62.700 72.800 ;
        RECT 58.000 72.100 58.600 72.200 ;
        RECT 58.200 71.100 58.600 72.100 ;
        RECT 59.700 71.800 60.200 72.200 ;
        RECT 59.800 71.100 60.200 71.800 ;
        RECT 63.000 71.100 63.400 73.100 ;
        RECT 65.400 71.100 65.800 73.100 ;
        RECT 66.200 73.000 68.200 73.100 ;
        RECT 66.200 71.100 66.600 73.000 ;
        RECT 67.800 71.100 68.200 73.000 ;
        RECT 72.000 71.100 72.400 73.900 ;
        RECT 73.400 71.100 73.800 74.800 ;
        RECT 75.100 74.200 75.400 75.800 ;
        RECT 76.200 74.800 77.000 75.200 ;
        RECT 77.400 75.100 77.800 76.200 ;
        RECT 78.200 75.900 80.200 76.200 ;
        RECT 80.600 75.900 81.000 79.900 ;
        RECT 81.400 76.900 81.800 79.900 ;
        RECT 81.500 76.600 81.800 76.900 ;
        RECT 83.000 79.600 85.000 79.900 ;
        RECT 83.000 76.900 83.400 79.600 ;
        RECT 83.800 76.900 84.200 79.300 ;
        RECT 84.600 77.000 85.000 79.600 ;
        RECT 85.500 79.600 87.300 79.900 ;
        RECT 85.500 79.500 85.800 79.600 ;
        RECT 83.000 76.600 83.300 76.900 ;
        RECT 81.500 76.300 83.300 76.600 ;
        RECT 83.900 76.700 84.200 76.900 ;
        RECT 85.400 76.700 85.800 79.500 ;
        RECT 87.000 79.500 87.300 79.600 ;
        RECT 83.900 76.500 85.800 76.700 ;
        RECT 86.200 76.500 86.600 79.300 ;
        RECT 87.000 76.500 87.400 79.500 ;
        RECT 83.900 76.400 85.700 76.500 ;
        RECT 86.200 76.200 86.500 76.500 ;
        RECT 87.800 76.200 88.200 79.900 ;
        RECT 90.200 76.200 90.600 79.900 ;
        RECT 92.600 76.200 93.000 79.900 ;
        RECT 96.600 76.200 97.000 79.900 ;
        RECT 86.200 76.100 86.600 76.200 ;
        RECT 78.600 75.200 79.000 75.400 ;
        RECT 80.600 75.200 80.900 75.900 ;
        RECT 84.900 75.800 86.600 76.100 ;
        RECT 87.800 75.900 88.900 76.200 ;
        RECT 90.200 75.900 91.300 76.200 ;
        RECT 92.600 75.900 93.700 76.200 ;
        RECT 78.200 75.100 79.000 75.200 ;
        RECT 77.400 74.900 79.000 75.100 ;
        RECT 79.800 74.900 81.000 75.200 ;
        RECT 77.400 74.800 78.600 74.900 ;
        RECT 75.100 74.100 75.900 74.200 ;
        RECT 75.100 73.900 76.000 74.100 ;
        RECT 74.200 72.400 74.600 73.200 ;
        RECT 75.600 72.100 76.000 73.900 ;
        RECT 79.000 73.800 79.400 74.600 ;
        RECT 79.800 74.100 80.100 74.900 ;
        RECT 80.600 74.800 81.000 74.900 ;
        RECT 83.800 74.800 84.600 75.200 ;
        RECT 84.900 75.100 85.200 75.800 ;
        RECT 88.600 75.600 88.900 75.900 ;
        RECT 91.000 75.600 91.300 75.900 ;
        RECT 93.400 75.600 93.700 75.900 ;
        RECT 95.900 75.900 97.000 76.200 ;
        RECT 95.900 75.600 96.200 75.900 ;
        RECT 88.600 75.200 89.200 75.600 ;
        RECT 91.000 75.200 91.600 75.600 ;
        RECT 93.400 75.200 94.000 75.600 ;
        RECT 95.600 75.200 96.200 75.600 ;
        RECT 87.800 75.100 88.200 75.200 ;
        RECT 84.900 74.800 88.200 75.100 ;
        RECT 83.000 74.100 83.800 74.200 ;
        RECT 79.800 73.800 83.800 74.100 ;
        RECT 76.600 72.800 77.000 73.200 ;
        RECT 79.800 73.100 80.100 73.800 ;
        RECT 80.600 73.100 81.000 73.200 ;
        RECT 81.400 73.100 81.800 73.200 ;
        RECT 76.600 72.100 76.900 72.800 ;
        RECT 75.600 71.800 76.900 72.100 ;
        RECT 75.600 71.100 76.000 71.800 ;
        RECT 79.800 71.100 80.200 73.100 ;
        RECT 80.600 72.800 81.800 73.100 ;
        RECT 82.200 72.800 83.100 73.200 ;
        RECT 80.500 72.400 80.900 72.800 ;
        RECT 84.900 72.500 85.200 74.800 ;
        RECT 87.800 74.400 88.200 74.800 ;
        RECT 88.600 73.700 88.900 75.200 ;
        RECT 90.200 74.400 90.600 75.200 ;
        RECT 91.000 73.700 91.300 75.200 ;
        RECT 92.600 74.400 93.000 75.200 ;
        RECT 93.400 73.700 93.700 75.200 ;
        RECT 83.200 72.200 85.200 72.500 ;
        RECT 83.200 72.100 83.500 72.200 ;
        RECT 83.000 71.800 83.500 72.100 ;
        RECT 84.600 72.100 85.200 72.200 ;
        RECT 87.800 73.400 88.900 73.700 ;
        RECT 90.200 73.400 91.300 73.700 ;
        RECT 92.600 73.400 93.700 73.700 ;
        RECT 95.900 73.700 96.200 75.200 ;
        RECT 96.600 74.400 97.000 75.200 ;
        RECT 95.900 73.400 97.000 73.700 ;
        RECT 83.000 71.100 83.400 71.800 ;
        RECT 84.600 71.100 85.000 72.100 ;
        RECT 87.800 71.100 88.200 73.400 ;
        RECT 90.200 71.100 90.600 73.400 ;
        RECT 92.600 71.100 93.000 73.400 ;
        RECT 96.600 71.100 97.000 73.400 ;
        RECT 3.000 68.900 3.400 69.900 ;
        RECT 4.600 69.200 5.000 69.900 ;
        RECT 2.800 68.800 3.400 68.900 ;
        RECT 4.500 68.800 5.000 69.200 ;
        RECT 2.800 68.500 4.800 68.800 ;
        RECT 2.800 65.200 3.100 68.500 ;
        RECT 7.300 68.200 7.700 69.900 ;
        RECT 10.200 68.900 10.600 69.900 ;
        RECT 4.900 67.800 5.800 68.200 ;
        RECT 7.300 67.900 8.200 68.200 ;
        RECT 4.200 66.800 5.000 67.200 ;
        RECT 3.400 65.800 4.200 66.200 ;
        RECT 7.800 66.100 8.200 67.900 ;
        RECT 8.600 67.100 9.000 67.600 ;
        RECT 10.200 67.200 10.500 68.900 ;
        RECT 11.000 67.800 11.400 68.600 ;
        RECT 12.400 67.200 12.800 69.900 ;
        RECT 15.300 68.200 15.700 69.900 ;
        RECT 17.700 68.200 18.100 69.900 ;
        RECT 20.600 68.900 21.000 69.900 ;
        RECT 15.300 67.900 16.200 68.200 ;
        RECT 17.700 67.900 18.600 68.200 ;
        RECT 10.200 67.100 10.600 67.200 ;
        RECT 8.600 66.800 10.600 67.100 ;
        RECT 11.800 66.900 12.800 67.200 ;
        RECT 11.800 66.800 12.700 66.900 ;
        RECT 7.800 65.800 8.900 66.100 ;
        RECT 1.400 64.900 3.100 65.200 ;
        RECT 1.400 64.800 1.800 64.900 ;
        RECT 1.500 64.500 1.800 64.800 ;
        RECT 2.300 64.500 4.100 64.600 ;
        RECT 0.600 61.500 1.000 64.500 ;
        RECT 1.400 61.700 1.800 64.500 ;
        RECT 2.200 64.300 4.100 64.500 ;
        RECT 0.700 61.400 1.000 61.500 ;
        RECT 2.200 61.500 2.600 64.300 ;
        RECT 3.800 64.100 4.100 64.300 ;
        RECT 4.700 64.400 6.500 64.700 ;
        RECT 7.000 64.400 7.400 65.200 ;
        RECT 4.700 64.100 5.000 64.400 ;
        RECT 2.200 61.400 2.500 61.500 ;
        RECT 0.700 61.100 2.500 61.400 ;
        RECT 3.000 61.400 3.400 64.000 ;
        RECT 3.800 61.700 4.200 64.100 ;
        RECT 4.600 61.400 5.000 64.100 ;
        RECT 3.000 61.100 5.000 61.400 ;
        RECT 6.200 64.100 6.500 64.400 ;
        RECT 6.200 61.100 6.600 64.100 ;
        RECT 7.800 61.100 8.200 65.800 ;
        RECT 8.600 65.200 8.900 65.800 ;
        RECT 9.400 65.400 9.800 66.200 ;
        RECT 8.600 64.800 9.000 65.200 ;
        RECT 10.200 65.100 10.500 66.800 ;
        RECT 11.900 65.200 12.200 66.800 ;
        RECT 13.000 65.800 13.800 66.200 ;
        RECT 9.700 64.700 10.600 65.100 ;
        RECT 11.800 64.800 12.200 65.200 ;
        RECT 14.200 64.800 14.600 65.600 ;
        RECT 9.700 61.100 10.100 64.700 ;
        RECT 11.900 63.500 12.200 64.800 ;
        RECT 12.600 63.800 13.000 64.600 ;
        RECT 15.000 64.400 15.400 65.200 ;
        RECT 11.900 63.200 13.700 63.500 ;
        RECT 11.900 63.100 12.200 63.200 ;
        RECT 11.800 61.100 12.200 63.100 ;
        RECT 13.400 63.100 13.700 63.200 ;
        RECT 13.400 61.100 13.800 63.100 ;
        RECT 15.800 61.100 16.200 67.900 ;
        RECT 16.600 66.800 17.000 67.600 ;
        RECT 17.400 66.800 17.800 67.200 ;
        RECT 17.400 66.100 17.700 66.800 ;
        RECT 18.200 66.100 18.600 67.900 ;
        RECT 19.800 67.800 20.200 68.600 ;
        RECT 20.700 67.200 21.000 68.900 ;
        RECT 20.600 66.800 21.000 67.200 ;
        RECT 17.400 65.800 18.600 66.100 ;
        RECT 17.400 64.400 17.800 65.200 ;
        RECT 18.200 61.100 18.600 65.800 ;
        RECT 20.700 65.100 21.000 66.800 ;
        RECT 23.000 68.900 23.400 69.900 ;
        RECT 25.400 68.900 25.800 69.900 ;
        RECT 29.400 68.900 29.800 69.900 ;
        RECT 31.800 68.900 32.200 69.900 ;
        RECT 34.200 68.900 34.600 69.900 ;
        RECT 36.600 68.900 37.000 69.900 ;
        RECT 23.000 67.200 23.300 68.900 ;
        RECT 23.800 67.800 24.200 68.600 ;
        RECT 24.600 67.800 25.000 68.600 ;
        RECT 25.500 67.200 25.800 68.900 ;
        RECT 28.600 67.800 29.000 68.600 ;
        RECT 29.500 67.200 29.800 68.900 ;
        RECT 30.200 68.100 30.600 68.200 ;
        RECT 31.000 68.100 31.400 68.600 ;
        RECT 30.200 67.800 31.400 68.100 ;
        RECT 31.900 67.200 32.200 68.900 ;
        RECT 32.600 68.100 33.000 68.200 ;
        RECT 33.400 68.100 33.800 68.600 ;
        RECT 32.600 67.800 33.800 68.100 ;
        RECT 34.300 67.200 34.600 68.900 ;
        RECT 35.800 67.800 36.200 68.600 ;
        RECT 36.700 67.200 37.000 68.900 ;
        RECT 23.000 66.800 23.400 67.200 ;
        RECT 25.400 66.800 25.800 67.200 ;
        RECT 29.400 66.800 29.800 67.200 ;
        RECT 31.800 66.800 32.200 67.200 ;
        RECT 34.200 66.800 34.600 67.200 ;
        RECT 36.600 66.800 37.000 67.200 ;
        RECT 21.400 66.100 21.800 66.200 ;
        RECT 22.200 66.100 22.600 66.200 ;
        RECT 21.400 65.800 22.600 66.100 ;
        RECT 21.400 65.400 21.800 65.800 ;
        RECT 22.200 65.400 22.600 65.800 ;
        RECT 23.000 66.100 23.300 66.800 ;
        RECT 23.800 66.100 24.200 66.200 ;
        RECT 23.000 65.800 24.200 66.100 ;
        RECT 23.000 65.100 23.300 65.800 ;
        RECT 25.500 65.100 25.800 66.800 ;
        RECT 26.200 65.400 26.600 66.200 ;
        RECT 29.500 65.200 29.800 66.800 ;
        RECT 30.200 65.400 30.600 66.200 ;
        RECT 29.400 65.100 29.800 65.200 ;
        RECT 31.900 65.100 32.200 66.800 ;
        RECT 32.600 65.400 33.000 66.200 ;
        RECT 34.300 65.100 34.600 66.800 ;
        RECT 35.000 65.400 35.400 66.200 ;
        RECT 36.700 65.100 37.000 66.800 ;
        RECT 39.000 68.900 39.400 69.900 ;
        RECT 41.400 68.900 41.800 69.900 ;
        RECT 39.000 67.200 39.300 68.900 ;
        RECT 39.800 67.800 40.200 68.600 ;
        RECT 41.500 67.200 41.800 68.900 ;
        RECT 39.000 66.800 39.400 67.200 ;
        RECT 41.400 66.800 41.800 67.200 ;
        RECT 43.000 66.800 43.400 67.600 ;
        RECT 37.400 66.100 37.800 66.200 ;
        RECT 38.200 66.100 38.600 66.200 ;
        RECT 37.400 65.800 38.600 66.100 ;
        RECT 37.400 65.400 37.800 65.800 ;
        RECT 38.200 65.400 38.600 65.800 ;
        RECT 39.000 65.100 39.300 66.800 ;
        RECT 41.500 65.100 41.800 66.800 ;
        RECT 42.200 65.400 42.600 66.200 ;
        RECT 20.600 64.700 21.500 65.100 ;
        RECT 21.100 62.200 21.500 64.700 ;
        RECT 22.500 64.700 23.400 65.100 ;
        RECT 25.400 64.700 26.300 65.100 ;
        RECT 29.400 64.700 30.300 65.100 ;
        RECT 31.800 64.700 32.700 65.100 ;
        RECT 34.200 64.700 35.100 65.100 ;
        RECT 36.600 64.700 37.500 65.100 ;
        RECT 22.500 64.200 22.900 64.700 ;
        RECT 22.200 63.800 22.900 64.200 ;
        RECT 21.100 61.800 21.800 62.200 ;
        RECT 21.100 61.100 21.500 61.800 ;
        RECT 22.500 61.100 22.900 63.800 ;
        RECT 25.900 62.200 26.300 64.700 ;
        RECT 25.900 61.800 26.600 62.200 ;
        RECT 25.900 61.100 26.300 61.800 ;
        RECT 29.900 61.100 30.300 64.700 ;
        RECT 32.300 62.200 32.700 64.700 ;
        RECT 34.700 62.200 35.100 64.700 ;
        RECT 37.100 62.200 37.500 64.700 ;
        RECT 38.500 64.700 39.400 65.100 ;
        RECT 41.400 64.700 42.300 65.100 ;
        RECT 38.500 64.200 38.900 64.700 ;
        RECT 38.200 63.800 38.900 64.200 ;
        RECT 32.300 61.800 33.000 62.200 ;
        RECT 34.700 61.800 35.400 62.200 ;
        RECT 37.100 61.800 37.800 62.200 ;
        RECT 32.300 61.100 32.700 61.800 ;
        RECT 34.700 61.100 35.100 61.800 ;
        RECT 37.100 61.100 37.500 61.800 ;
        RECT 38.500 61.100 38.900 63.800 ;
        RECT 41.900 62.200 42.300 64.700 ;
        RECT 41.400 61.800 42.300 62.200 ;
        RECT 41.900 61.100 42.300 61.800 ;
        RECT 43.800 61.100 44.200 69.900 ;
        RECT 45.900 67.900 46.700 69.900 ;
        RECT 48.600 67.900 49.000 69.900 ;
        RECT 49.400 68.000 49.800 69.900 ;
        RECT 51.000 68.000 51.400 69.900 ;
        RECT 49.400 67.900 51.400 68.000 ;
        RECT 45.400 66.800 45.800 67.200 ;
        RECT 45.500 66.600 45.800 66.800 ;
        RECT 45.500 66.200 45.900 66.600 ;
        RECT 46.200 66.200 46.500 67.900 ;
        RECT 48.700 67.200 49.000 67.900 ;
        RECT 49.500 67.700 51.300 67.900 ;
        RECT 50.600 67.200 51.000 67.400 ;
        RECT 47.000 66.400 47.400 67.200 ;
        RECT 48.600 66.800 49.900 67.200 ;
        RECT 50.600 66.900 51.400 67.200 ;
        RECT 51.000 66.800 51.400 66.900 ;
        RECT 51.800 66.800 52.200 67.600 ;
        RECT 52.600 67.100 53.000 69.900 ;
        RECT 53.500 68.200 53.900 68.600 ;
        RECT 53.400 67.800 53.800 68.200 ;
        RECT 54.200 67.900 54.600 69.900 ;
        RECT 56.600 67.900 57.000 69.900 ;
        RECT 57.400 68.000 57.800 69.900 ;
        RECT 59.000 68.000 59.400 69.900 ;
        RECT 57.400 67.900 59.400 68.000 ;
        RECT 59.800 68.000 60.200 69.900 ;
        RECT 61.400 69.600 63.400 69.900 ;
        RECT 61.400 68.000 61.800 69.600 ;
        RECT 59.800 67.900 61.800 68.000 ;
        RECT 53.400 67.100 53.800 67.200 ;
        RECT 52.600 66.800 53.800 67.100 ;
        RECT 44.600 65.400 45.000 66.200 ;
        RECT 46.200 65.800 46.600 66.200 ;
        RECT 47.800 66.100 48.200 66.200 ;
        RECT 47.400 65.800 48.200 66.100 ;
        RECT 46.200 65.700 46.500 65.800 ;
        RECT 45.500 65.400 46.500 65.700 ;
        RECT 47.400 65.600 47.800 65.800 ;
        RECT 45.500 65.100 45.800 65.400 ;
        RECT 49.600 65.200 49.900 66.800 ;
        RECT 50.200 65.800 50.600 66.600 ;
        RECT 48.600 65.100 49.000 65.200 ;
        RECT 44.600 61.400 45.000 65.100 ;
        RECT 45.400 61.700 45.800 65.100 ;
        RECT 46.200 64.800 48.200 65.100 ;
        RECT 48.600 64.800 49.300 65.100 ;
        RECT 49.600 64.800 50.600 65.200 ;
        RECT 46.200 61.400 46.600 64.800 ;
        RECT 44.600 61.100 46.600 61.400 ;
        RECT 47.800 61.100 48.200 64.800 ;
        RECT 49.000 64.200 49.300 64.800 ;
        RECT 49.000 63.800 49.400 64.200 ;
        RECT 49.700 61.100 50.100 64.800 ;
        RECT 52.600 61.100 53.000 66.800 ;
        RECT 53.400 66.100 53.800 66.200 ;
        RECT 54.300 66.100 54.600 67.900 ;
        RECT 56.700 67.200 57.000 67.900 ;
        RECT 57.500 67.700 59.300 67.900 ;
        RECT 59.900 67.700 61.700 67.900 ;
        RECT 62.200 67.800 62.600 69.300 ;
        RECT 63.000 67.900 63.400 69.600 ;
        RECT 64.600 68.900 65.000 69.900 ;
        RECT 63.800 67.800 64.200 68.600 ;
        RECT 58.600 67.200 59.000 67.400 ;
        RECT 60.200 67.200 60.600 67.400 ;
        RECT 62.300 67.200 62.600 67.800 ;
        RECT 64.700 67.200 65.000 68.900 ;
        RECT 55.000 66.400 55.400 67.200 ;
        RECT 56.600 66.800 57.900 67.200 ;
        RECT 58.600 66.900 59.400 67.200 ;
        RECT 59.000 66.800 59.400 66.900 ;
        RECT 59.800 66.900 60.600 67.200 ;
        RECT 61.400 66.900 62.600 67.200 ;
        RECT 59.800 66.800 60.200 66.900 ;
        RECT 61.400 66.800 61.800 66.900 ;
        RECT 55.800 66.100 56.200 66.200 ;
        RECT 53.400 65.800 54.600 66.100 ;
        RECT 55.400 65.800 56.200 66.100 ;
        RECT 53.500 65.100 53.800 65.800 ;
        RECT 55.400 65.600 55.800 65.800 ;
        RECT 56.600 65.100 57.000 65.200 ;
        RECT 57.600 65.100 57.900 66.800 ;
        RECT 58.200 66.100 58.600 66.600 ;
        RECT 59.000 66.100 59.400 66.200 ;
        RECT 58.200 65.800 59.400 66.100 ;
        RECT 60.600 65.800 61.000 66.600 ;
        RECT 61.400 65.100 61.700 66.800 ;
        RECT 62.200 65.800 62.600 66.600 ;
        RECT 63.000 66.400 63.400 67.200 ;
        RECT 64.600 66.800 65.000 67.200 ;
        RECT 66.200 66.800 66.600 67.600 ;
        RECT 64.700 65.100 65.000 66.800 ;
        RECT 65.400 65.400 65.800 66.200 ;
        RECT 53.400 61.100 53.800 65.100 ;
        RECT 54.200 64.800 56.200 65.100 ;
        RECT 56.600 64.800 57.300 65.100 ;
        RECT 57.600 64.800 58.100 65.100 ;
        RECT 54.200 61.100 54.600 64.800 ;
        RECT 55.800 61.100 56.200 64.800 ;
        RECT 57.000 64.200 57.300 64.800 ;
        RECT 57.000 63.800 57.400 64.200 ;
        RECT 57.700 62.200 58.100 64.800 ;
        RECT 57.700 61.800 58.600 62.200 ;
        RECT 57.700 61.100 58.100 61.800 ;
        RECT 61.100 61.100 62.100 65.100 ;
        RECT 64.600 64.700 65.500 65.100 ;
        RECT 65.100 64.200 65.500 64.700 ;
        RECT 65.100 63.800 65.800 64.200 ;
        RECT 65.100 61.100 65.500 63.800 ;
        RECT 67.000 62.100 67.400 69.900 ;
        RECT 71.200 67.100 71.600 69.900 ;
        RECT 73.900 69.200 74.300 69.900 ;
        RECT 73.400 68.800 74.300 69.200 ;
        RECT 73.900 68.200 74.300 68.800 ;
        RECT 73.400 67.900 74.300 68.200 ;
        RECT 75.000 68.000 75.400 69.900 ;
        RECT 76.600 68.000 77.000 69.900 ;
        RECT 75.000 67.900 77.000 68.000 ;
        RECT 77.400 67.900 77.800 69.900 ;
        RECT 79.000 68.900 79.400 69.900 ;
        RECT 71.200 66.900 72.100 67.100 ;
        RECT 71.300 66.800 72.100 66.900 ;
        RECT 72.600 66.800 73.000 67.600 ;
        RECT 70.200 65.800 71.400 66.200 ;
        RECT 68.600 65.100 69.000 65.200 ;
        RECT 69.400 65.100 69.800 65.600 ;
        RECT 68.600 64.800 69.800 65.100 ;
        RECT 71.800 65.200 72.100 66.800 ;
        RECT 71.800 64.800 72.200 65.200 ;
        RECT 71.000 63.800 71.400 64.600 ;
        RECT 71.800 63.500 72.100 64.800 ;
        RECT 70.300 63.200 72.100 63.500 ;
        RECT 68.600 62.100 69.000 62.200 ;
        RECT 67.000 61.800 69.000 62.100 ;
        RECT 67.000 61.100 67.400 61.800 ;
        RECT 70.200 61.100 70.600 63.200 ;
        RECT 71.800 63.100 72.100 63.200 ;
        RECT 71.800 61.100 72.200 63.100 ;
        RECT 73.400 61.100 73.800 67.900 ;
        RECT 75.100 67.700 76.900 67.900 ;
        RECT 75.400 67.200 75.800 67.400 ;
        RECT 77.400 67.200 77.700 67.900 ;
        RECT 79.100 67.200 79.400 68.900 ;
        RECT 81.400 68.800 81.800 69.900 ;
        RECT 80.600 67.800 81.000 68.600 ;
        RECT 81.500 67.200 81.800 68.800 ;
        RECT 75.000 66.900 75.800 67.200 ;
        RECT 75.000 66.800 75.400 66.900 ;
        RECT 76.500 66.800 77.800 67.200 ;
        RECT 78.200 67.100 78.600 67.200 ;
        RECT 79.000 67.100 79.400 67.200 ;
        RECT 78.200 66.800 79.400 67.100 ;
        RECT 81.400 66.800 81.800 67.200 ;
        RECT 83.600 67.100 84.000 69.900 ;
        RECT 86.300 68.200 86.700 68.600 ;
        RECT 86.200 67.800 86.600 68.200 ;
        RECT 87.000 67.900 87.400 69.900 ;
        RECT 89.500 68.200 89.900 68.600 ;
        RECT 74.200 66.100 74.600 66.200 ;
        RECT 75.800 66.100 76.200 66.600 ;
        RECT 74.200 65.800 76.200 66.100 ;
        RECT 74.200 64.400 74.600 65.200 ;
        RECT 76.500 65.100 76.800 66.800 ;
        RECT 77.400 65.100 77.800 65.200 ;
        RECT 79.100 65.100 79.400 66.800 ;
        RECT 79.800 65.400 80.200 66.200 ;
        RECT 80.600 66.100 81.000 66.200 ;
        RECT 81.500 66.100 81.800 66.800 ;
        RECT 83.100 66.900 84.000 67.100 ;
        RECT 86.200 67.100 86.600 67.200 ;
        RECT 87.100 67.100 87.400 67.900 ;
        RECT 89.400 67.800 89.800 68.200 ;
        RECT 90.200 67.900 90.600 69.900 ;
        RECT 83.100 66.800 83.900 66.900 ;
        RECT 86.200 66.800 87.400 67.100 ;
        RECT 80.600 65.800 81.800 66.100 ;
        RECT 81.500 65.100 81.800 65.800 ;
        RECT 82.200 65.400 82.600 66.200 ;
        RECT 83.100 65.200 83.400 66.800 ;
        RECT 84.200 65.800 85.000 66.200 ;
        RECT 86.200 66.100 86.600 66.200 ;
        RECT 87.100 66.100 87.400 66.800 ;
        RECT 87.800 66.400 88.200 67.200 ;
        RECT 88.600 66.100 89.000 66.200 ;
        RECT 86.200 65.800 87.400 66.100 ;
        RECT 88.200 65.800 89.000 66.100 ;
        RECT 89.400 66.100 89.800 66.200 ;
        RECT 90.300 66.100 90.600 67.900 ;
        RECT 91.000 66.400 91.400 67.200 ;
        RECT 91.800 66.100 92.200 66.200 ;
        RECT 89.400 65.800 90.600 66.100 ;
        RECT 91.400 65.800 92.200 66.100 ;
        RECT 76.300 64.800 76.800 65.100 ;
        RECT 77.100 64.800 77.800 65.100 ;
        RECT 76.300 64.200 76.700 64.800 ;
        RECT 77.100 64.200 77.400 64.800 ;
        RECT 79.000 64.700 79.900 65.100 ;
        RECT 81.400 64.700 82.300 65.100 ;
        RECT 83.000 64.800 83.400 65.200 ;
        RECT 85.400 64.800 85.800 65.600 ;
        RECT 86.300 65.100 86.600 65.800 ;
        RECT 88.200 65.600 88.600 65.800 ;
        RECT 89.500 65.100 89.800 65.800 ;
        RECT 91.400 65.600 91.800 65.800 ;
        RECT 75.800 63.800 76.700 64.200 ;
        RECT 77.000 63.800 77.400 64.200 ;
        RECT 76.300 61.100 76.700 63.800 ;
        RECT 79.500 61.100 79.900 64.700 ;
        RECT 81.900 61.100 82.300 64.700 ;
        RECT 83.100 63.500 83.400 64.800 ;
        RECT 83.800 63.800 84.200 64.600 ;
        RECT 83.100 63.200 84.900 63.500 ;
        RECT 83.100 63.100 83.400 63.200 ;
        RECT 83.000 61.100 83.400 63.100 ;
        RECT 84.600 61.100 85.000 63.200 ;
        RECT 86.200 61.100 86.600 65.100 ;
        RECT 87.000 64.800 89.000 65.100 ;
        RECT 87.000 61.100 87.400 64.800 ;
        RECT 88.600 61.100 89.000 64.800 ;
        RECT 89.400 61.100 89.800 65.100 ;
        RECT 90.200 64.800 92.200 65.100 ;
        RECT 90.200 61.100 90.600 64.800 ;
        RECT 91.800 61.100 92.200 64.800 ;
        RECT 92.600 61.100 93.000 69.900 ;
        RECT 93.400 67.800 93.800 68.600 ;
        RECT 94.500 68.200 94.900 69.900 ;
        RECT 94.500 67.900 95.400 68.200 ;
        RECT 95.000 66.100 95.400 67.900 ;
        RECT 95.800 66.800 96.200 67.600 ;
        RECT 96.600 66.100 97.000 66.200 ;
        RECT 95.000 65.800 97.000 66.100 ;
        RECT 94.200 64.400 94.600 65.200 ;
        RECT 95.000 61.100 95.400 65.800 ;
        RECT 1.400 55.100 1.800 59.900 ;
        RECT 3.800 57.900 4.200 59.900 ;
        RECT 3.900 57.800 4.200 57.900 ;
        RECT 5.400 57.900 5.800 59.900 ;
        RECT 7.000 57.900 7.400 59.900 ;
        RECT 5.400 57.800 5.700 57.900 ;
        RECT 3.900 57.500 5.700 57.800 ;
        RECT 2.200 55.800 2.600 56.600 ;
        RECT 4.600 56.400 5.000 57.200 ;
        RECT 5.400 56.200 5.700 57.500 ;
        RECT 3.000 55.100 3.400 56.200 ;
        RECT 5.400 55.800 5.800 56.200 ;
        RECT 7.100 55.800 7.400 57.900 ;
        RECT 8.600 55.900 9.000 59.900 ;
        RECT 10.700 55.900 11.700 59.900 ;
        RECT 1.400 54.800 3.400 55.100 ;
        RECT 3.800 54.800 4.600 55.200 ;
        RECT 1.400 53.100 1.800 54.800 ;
        RECT 5.400 54.200 5.700 55.800 ;
        RECT 7.100 55.500 8.300 55.800 ;
        RECT 4.900 54.100 5.700 54.200 ;
        RECT 4.800 53.900 5.700 54.100 ;
        RECT 1.400 52.800 2.300 53.100 ;
        RECT 1.900 51.100 2.300 52.800 ;
        RECT 4.800 51.100 5.200 53.900 ;
        RECT 8.000 53.800 8.300 55.500 ;
        RECT 8.700 55.200 9.000 55.900 ;
        RECT 8.600 54.800 9.000 55.200 ;
        RECT 8.000 53.700 8.400 53.800 ;
        RECT 6.900 53.500 8.400 53.700 ;
        RECT 6.300 53.400 8.400 53.500 ;
        RECT 6.300 53.200 7.200 53.400 ;
        RECT 6.300 53.100 6.600 53.200 ;
        RECT 8.700 53.100 9.000 54.800 ;
        RECT 9.400 53.800 9.800 54.600 ;
        RECT 10.200 54.400 10.600 55.200 ;
        RECT 11.100 54.200 11.400 55.900 ;
        RECT 11.800 54.400 12.200 55.200 ;
        RECT 11.000 54.100 11.400 54.200 ;
        RECT 10.200 53.800 11.400 54.100 ;
        RECT 10.200 53.100 10.500 53.800 ;
        RECT 11.100 53.100 12.900 53.300 ;
        RECT 14.200 53.100 14.600 59.900 ;
        RECT 6.200 51.100 6.600 53.100 ;
        RECT 8.300 52.600 9.000 53.100 ;
        RECT 8.300 52.200 8.700 52.600 ;
        RECT 8.300 51.800 9.000 52.200 ;
        RECT 8.300 51.100 8.700 51.800 ;
        RECT 9.400 51.400 9.800 53.100 ;
        RECT 10.200 51.700 10.600 53.100 ;
        RECT 11.000 53.000 13.000 53.100 ;
        RECT 11.000 51.400 11.400 53.000 ;
        RECT 9.400 51.100 11.400 51.400 ;
        RECT 12.600 51.100 13.000 53.000 ;
        RECT 14.200 52.800 15.100 53.100 ;
        RECT 14.700 51.100 15.100 52.800 ;
        RECT 16.600 51.100 17.000 59.900 ;
        RECT 18.700 56.200 19.100 59.900 ;
        RECT 21.400 57.900 21.800 59.900 ;
        RECT 21.500 57.800 21.800 57.900 ;
        RECT 23.000 57.900 23.400 59.900 ;
        RECT 24.900 59.200 25.300 59.900 ;
        RECT 24.900 58.800 25.800 59.200 ;
        RECT 23.000 57.800 23.300 57.900 ;
        RECT 21.500 57.500 23.300 57.800 ;
        RECT 19.400 56.800 19.800 57.200 ;
        RECT 19.500 56.200 19.800 56.800 ;
        RECT 22.200 56.400 22.600 57.200 ;
        RECT 23.000 56.200 23.300 57.500 ;
        RECT 24.200 56.800 24.600 57.200 ;
        RECT 24.200 56.200 24.500 56.800 ;
        RECT 24.900 56.200 25.300 58.800 ;
        RECT 18.700 55.900 19.200 56.200 ;
        RECT 19.500 55.900 20.200 56.200 ;
        RECT 18.200 54.400 18.600 55.200 ;
        RECT 18.900 55.100 19.200 55.900 ;
        RECT 19.800 55.800 20.200 55.900 ;
        RECT 20.600 55.100 21.000 56.200 ;
        RECT 23.000 56.100 23.400 56.200 ;
        RECT 23.800 56.100 24.500 56.200 ;
        RECT 23.000 55.900 24.500 56.100 ;
        RECT 24.800 55.900 25.300 56.200 ;
        RECT 28.900 56.300 29.300 59.900 ;
        RECT 28.900 55.900 29.800 56.300 ;
        RECT 23.000 55.800 24.200 55.900 ;
        RECT 18.900 54.800 21.000 55.100 ;
        RECT 21.400 54.800 22.200 55.200 ;
        RECT 18.900 54.200 19.200 54.800 ;
        RECT 23.000 54.200 23.300 55.800 ;
        RECT 24.800 54.200 25.100 55.900 ;
        RECT 25.400 55.100 25.800 55.200 ;
        RECT 25.400 54.800 27.300 55.100 ;
        RECT 28.600 54.800 29.000 55.600 ;
        RECT 25.400 54.400 25.800 54.800 ;
        RECT 17.400 54.100 17.800 54.200 ;
        RECT 17.400 53.800 18.200 54.100 ;
        RECT 18.900 53.800 20.200 54.200 ;
        RECT 22.500 54.100 23.300 54.200 ;
        RECT 22.400 53.900 23.300 54.100 ;
        RECT 17.800 53.600 18.200 53.800 ;
        RECT 17.500 53.100 19.300 53.300 ;
        RECT 19.800 53.100 20.100 53.800 ;
        RECT 17.400 53.000 19.400 53.100 ;
        RECT 17.400 51.100 17.800 53.000 ;
        RECT 19.000 51.100 19.400 53.000 ;
        RECT 19.800 51.100 20.200 53.100 ;
        RECT 22.400 51.100 22.800 53.900 ;
        RECT 23.800 53.800 25.100 54.200 ;
        RECT 26.200 54.100 26.600 54.200 ;
        RECT 25.800 53.800 26.600 54.100 ;
        RECT 27.000 54.100 27.300 54.800 ;
        RECT 29.400 54.200 29.700 55.900 ;
        RECT 31.000 55.800 31.400 56.600 ;
        RECT 29.400 54.100 29.800 54.200 ;
        RECT 27.000 53.800 29.800 54.100 ;
        RECT 23.900 53.100 24.200 53.800 ;
        RECT 25.800 53.600 26.200 53.800 ;
        RECT 24.700 53.100 26.500 53.300 ;
        RECT 23.800 51.100 24.200 53.100 ;
        RECT 24.600 53.000 26.600 53.100 ;
        RECT 24.600 51.100 25.000 53.000 ;
        RECT 26.200 51.100 26.600 53.000 ;
        RECT 29.400 52.100 29.700 53.800 ;
        RECT 30.200 53.100 30.600 53.200 ;
        RECT 31.800 53.100 32.200 59.900 ;
        RECT 30.200 52.800 32.200 53.100 ;
        RECT 34.200 54.100 34.600 59.900 ;
        RECT 35.000 56.200 35.400 59.900 ;
        RECT 36.600 59.600 38.600 59.900 ;
        RECT 36.600 56.200 37.000 59.600 ;
        RECT 35.000 55.900 37.000 56.200 ;
        RECT 37.400 55.900 37.800 59.300 ;
        RECT 38.200 55.900 38.600 59.600 ;
        RECT 39.400 56.800 39.800 57.200 ;
        RECT 39.400 56.200 39.700 56.800 ;
        RECT 40.100 56.200 40.500 59.900 ;
        RECT 39.000 55.900 39.700 56.200 ;
        RECT 40.000 55.900 40.500 56.200 ;
        RECT 42.500 56.300 42.900 59.900 ;
        RECT 45.000 56.800 45.400 57.200 ;
        RECT 42.500 55.900 43.400 56.300 ;
        RECT 45.000 56.200 45.300 56.800 ;
        RECT 45.700 56.200 46.100 59.900 ;
        RECT 44.600 55.900 45.300 56.200 ;
        RECT 45.600 55.900 46.100 56.200 ;
        RECT 37.400 55.600 37.700 55.900 ;
        RECT 39.000 55.800 39.400 55.900 ;
        RECT 35.400 55.200 35.800 55.400 ;
        RECT 36.700 55.300 37.700 55.600 ;
        RECT 36.700 55.200 37.000 55.300 ;
        RECT 35.000 54.900 35.800 55.200 ;
        RECT 35.000 54.800 35.400 54.900 ;
        RECT 36.600 54.800 37.000 55.200 ;
        RECT 38.200 55.100 38.600 55.600 ;
        RECT 40.000 55.100 40.300 55.900 ;
        RECT 38.200 54.800 40.300 55.100 ;
        RECT 35.800 54.100 36.200 54.600 ;
        RECT 34.200 53.800 36.200 54.100 ;
        RECT 30.200 52.400 30.600 52.800 ;
        RECT 29.400 51.100 29.800 52.100 ;
        RECT 31.300 51.100 31.700 52.800 ;
        RECT 34.200 51.100 34.600 53.800 ;
        RECT 36.700 53.100 37.000 54.800 ;
        RECT 37.300 54.400 37.700 54.800 ;
        RECT 37.400 54.200 37.700 54.400 ;
        RECT 40.000 54.200 40.300 54.800 ;
        RECT 40.600 55.100 41.000 55.200 ;
        RECT 41.400 55.100 41.800 55.200 ;
        RECT 40.600 54.800 41.800 55.100 ;
        RECT 42.200 54.800 42.600 55.600 ;
        RECT 43.000 55.100 43.300 55.900 ;
        RECT 44.600 55.800 45.000 55.900 ;
        RECT 44.600 55.100 44.900 55.800 ;
        RECT 43.000 54.800 44.900 55.100 ;
        RECT 40.600 54.400 41.000 54.800 ;
        RECT 43.000 54.200 43.300 54.800 ;
        RECT 45.600 54.200 45.900 55.900 ;
        RECT 46.200 54.400 46.600 55.200 ;
        RECT 37.400 53.800 37.800 54.200 ;
        RECT 39.000 53.800 40.300 54.200 ;
        RECT 41.400 54.100 41.800 54.200 ;
        RECT 41.000 53.800 41.800 54.100 ;
        RECT 43.000 53.800 43.400 54.200 ;
        RECT 44.600 53.800 45.900 54.200 ;
        RECT 47.000 54.100 47.400 54.200 ;
        RECT 46.600 53.800 47.400 54.100 ;
        RECT 39.100 53.100 39.400 53.800 ;
        RECT 41.000 53.600 41.400 53.800 ;
        RECT 39.900 53.100 41.700 53.300 ;
        RECT 36.500 51.100 37.300 53.100 ;
        RECT 39.000 51.100 39.400 53.100 ;
        RECT 39.800 53.000 41.800 53.100 ;
        RECT 39.800 51.100 40.200 53.000 ;
        RECT 41.400 51.100 41.800 53.000 ;
        RECT 43.000 52.100 43.300 53.800 ;
        RECT 43.800 52.400 44.200 53.200 ;
        RECT 44.700 53.100 45.000 53.800 ;
        RECT 46.600 53.600 47.000 53.800 ;
        RECT 45.500 53.100 47.300 53.300 ;
        RECT 43.000 51.100 43.400 52.100 ;
        RECT 44.600 51.100 45.000 53.100 ;
        RECT 45.400 53.000 47.400 53.100 ;
        RECT 45.400 51.100 45.800 53.000 ;
        RECT 47.000 51.100 47.400 53.000 ;
        RECT 47.800 52.400 48.200 53.200 ;
        RECT 48.600 51.100 49.000 59.900 ;
        RECT 49.400 55.800 49.800 56.600 ;
        RECT 50.200 53.100 50.600 59.900 ;
        RECT 52.200 56.800 52.600 57.200 ;
        RECT 52.200 56.200 52.500 56.800 ;
        RECT 52.900 56.200 53.300 59.900 ;
        RECT 55.400 56.800 55.800 57.200 ;
        RECT 55.400 56.200 55.700 56.800 ;
        RECT 56.100 56.200 56.500 59.900 ;
        RECT 51.800 55.900 52.500 56.200 ;
        RECT 52.800 55.900 53.300 56.200 ;
        RECT 55.000 55.900 55.700 56.200 ;
        RECT 56.000 55.900 56.500 56.200 ;
        RECT 58.500 56.300 58.900 59.900 ;
        RECT 58.500 55.900 59.400 56.300 ;
        RECT 61.900 55.900 62.900 59.900 ;
        RECT 64.600 57.100 65.000 59.900 ;
        RECT 64.600 56.800 65.700 57.100 ;
        RECT 51.800 55.800 52.200 55.900 ;
        RECT 51.800 55.100 52.200 55.200 ;
        RECT 52.800 55.100 53.100 55.900 ;
        RECT 55.000 55.800 55.400 55.900 ;
        RECT 51.800 54.800 53.100 55.100 ;
        RECT 52.800 54.200 53.100 54.800 ;
        RECT 53.400 54.400 53.800 55.200 ;
        RECT 56.000 54.200 56.300 55.900 ;
        RECT 56.600 54.400 57.000 55.200 ;
        RECT 58.200 54.800 58.600 55.600 ;
        RECT 59.000 54.200 59.300 55.900 ;
        RECT 59.800 54.800 61.000 55.100 ;
        RECT 59.800 54.200 60.100 54.800 ;
        RECT 51.000 53.400 51.400 54.200 ;
        RECT 51.800 53.800 53.100 54.200 ;
        RECT 54.200 54.100 54.600 54.200 ;
        RECT 55.000 54.100 56.300 54.200 ;
        RECT 57.400 54.100 57.800 54.200 ;
        RECT 58.200 54.100 58.600 54.200 ;
        RECT 53.800 53.800 56.300 54.100 ;
        RECT 57.000 53.800 58.600 54.100 ;
        RECT 59.000 53.800 59.400 54.200 ;
        RECT 59.800 53.800 60.200 54.200 ;
        RECT 60.600 53.800 61.000 54.800 ;
        RECT 61.400 54.400 61.800 55.200 ;
        RECT 62.300 54.200 62.600 55.900 ;
        RECT 63.000 55.100 63.400 55.200 ;
        RECT 64.600 55.100 65.000 56.800 ;
        RECT 65.400 56.200 65.700 56.800 ;
        RECT 67.500 56.300 67.900 59.900 ;
        RECT 65.400 55.800 65.800 56.200 ;
        RECT 67.000 55.900 67.900 56.300 ;
        RECT 70.500 56.300 70.900 59.900 ;
        RECT 73.400 57.900 73.800 59.900 ;
        RECT 73.500 57.800 73.800 57.900 ;
        RECT 75.000 57.900 75.400 59.900 ;
        RECT 75.000 57.800 75.300 57.900 ;
        RECT 73.500 57.500 75.300 57.800 ;
        RECT 74.200 56.400 74.600 57.200 ;
        RECT 70.500 55.900 71.400 56.300 ;
        RECT 75.000 56.200 75.300 57.500 ;
        RECT 77.100 56.300 77.500 59.900 ;
        RECT 79.500 56.300 79.900 59.900 ;
        RECT 63.000 54.800 65.000 55.100 ;
        RECT 63.000 54.400 63.400 54.800 ;
        RECT 62.200 54.100 62.600 54.200 ;
        RECT 63.800 54.100 64.200 54.200 ;
        RECT 61.400 53.800 62.600 54.100 ;
        RECT 63.400 53.800 64.200 54.100 ;
        RECT 51.900 53.100 52.200 53.800 ;
        RECT 53.800 53.600 54.200 53.800 ;
        RECT 52.700 53.100 54.500 53.300 ;
        RECT 55.100 53.100 55.400 53.800 ;
        RECT 57.000 53.600 57.400 53.800 ;
        RECT 55.900 53.100 57.700 53.300 ;
        RECT 49.700 52.800 50.600 53.100 ;
        RECT 49.700 51.100 50.100 52.800 ;
        RECT 51.800 51.100 52.200 53.100 ;
        RECT 52.600 53.000 54.600 53.100 ;
        RECT 52.600 51.100 53.000 53.000 ;
        RECT 54.200 51.100 54.600 53.000 ;
        RECT 55.000 51.100 55.400 53.100 ;
        RECT 55.800 53.000 57.800 53.100 ;
        RECT 55.800 51.100 56.200 53.000 ;
        RECT 57.400 51.100 57.800 53.000 ;
        RECT 59.000 52.200 59.300 53.800 ;
        RECT 61.400 53.200 61.700 53.800 ;
        RECT 63.400 53.600 63.800 53.800 ;
        RECT 59.800 52.400 60.200 53.200 ;
        RECT 59.000 51.100 59.400 52.200 ;
        RECT 60.600 51.400 61.000 53.100 ;
        RECT 61.400 51.700 61.800 53.200 ;
        RECT 62.300 53.100 64.100 53.300 ;
        RECT 62.200 53.000 64.200 53.100 ;
        RECT 62.200 51.400 62.600 53.000 ;
        RECT 60.600 51.100 62.600 51.400 ;
        RECT 63.800 51.100 64.200 53.000 ;
        RECT 64.600 51.100 65.000 54.800 ;
        RECT 67.100 54.200 67.400 55.900 ;
        RECT 67.800 55.100 68.200 55.600 ;
        RECT 69.400 55.100 69.800 55.200 ;
        RECT 67.800 54.800 69.800 55.100 ;
        RECT 70.200 54.800 70.600 55.600 ;
        RECT 67.000 53.800 67.400 54.200 ;
        RECT 65.400 52.400 65.800 53.200 ;
        RECT 66.200 52.400 66.600 53.200 ;
        RECT 67.100 52.200 67.400 53.800 ;
        RECT 67.000 51.100 67.400 52.200 ;
        RECT 71.000 54.200 71.300 55.900 ;
        RECT 72.600 55.400 73.000 56.200 ;
        RECT 75.000 55.800 75.400 56.200 ;
        RECT 76.600 55.900 77.500 56.300 ;
        RECT 79.000 55.900 79.900 56.300 ;
        RECT 81.000 56.800 81.400 57.200 ;
        RECT 81.000 56.200 81.300 56.800 ;
        RECT 81.700 56.200 82.100 59.900 ;
        RECT 80.600 55.900 81.300 56.200 ;
        RECT 81.600 55.900 82.100 56.200 ;
        RECT 84.100 56.300 84.500 59.900 ;
        RECT 87.300 59.200 87.700 59.900 ;
        RECT 87.300 58.800 88.200 59.200 ;
        RECT 86.600 56.800 87.000 57.200 ;
        RECT 84.100 55.900 85.000 56.300 ;
        RECT 86.600 56.200 86.900 56.800 ;
        RECT 87.300 56.200 87.700 58.800 ;
        RECT 73.400 54.800 74.200 55.200 ;
        RECT 75.000 54.200 75.300 55.800 ;
        RECT 71.000 53.800 71.400 54.200 ;
        RECT 74.500 54.100 75.300 54.200 ;
        RECT 74.400 53.900 75.300 54.100 ;
        RECT 75.800 54.800 76.200 55.200 ;
        RECT 75.800 54.100 76.100 54.800 ;
        RECT 76.700 54.200 77.000 55.900 ;
        RECT 77.400 54.800 77.800 55.600 ;
        RECT 79.100 55.200 79.400 55.900 ;
        RECT 80.600 55.800 81.000 55.900 ;
        RECT 81.600 55.200 81.900 55.900 ;
        RECT 84.600 55.800 85.000 55.900 ;
        RECT 86.200 55.900 86.900 56.200 ;
        RECT 87.200 55.900 87.700 56.200 ;
        RECT 86.200 55.800 86.600 55.900 ;
        RECT 79.000 54.800 79.400 55.200 ;
        RECT 81.400 54.800 81.900 55.200 ;
        RECT 79.100 54.200 79.400 54.800 ;
        RECT 81.600 54.200 81.900 54.800 ;
        RECT 82.200 54.400 82.600 55.200 ;
        RECT 83.000 55.100 83.400 55.200 ;
        RECT 83.800 55.100 84.200 55.600 ;
        RECT 83.000 54.800 84.200 55.100 ;
        RECT 84.600 54.200 84.900 55.800 ;
        RECT 87.200 54.200 87.500 55.900 ;
        RECT 87.800 54.400 88.200 55.200 ;
        RECT 76.600 54.100 77.000 54.200 ;
        RECT 71.000 53.200 71.300 53.800 ;
        RECT 71.000 52.800 71.400 53.200 ;
        RECT 71.000 52.100 71.300 52.800 ;
        RECT 71.800 52.400 72.200 53.200 ;
        RECT 71.000 51.100 71.400 52.100 ;
        RECT 74.400 51.100 74.800 53.900 ;
        RECT 75.800 53.800 77.000 54.100 ;
        RECT 79.000 53.800 79.400 54.200 ;
        RECT 80.600 53.800 81.900 54.200 ;
        RECT 83.000 54.100 83.400 54.200 ;
        RECT 82.600 53.800 83.400 54.100 ;
        RECT 84.600 53.800 85.000 54.200 ;
        RECT 86.200 53.800 87.500 54.200 ;
        RECT 88.600 54.100 89.000 54.200 ;
        RECT 89.400 54.100 89.800 59.900 ;
        RECT 88.200 53.800 89.800 54.100 ;
        RECT 75.800 52.400 76.200 53.200 ;
        RECT 76.700 52.100 77.000 53.800 ;
        RECT 79.100 52.100 79.400 53.800 ;
        RECT 80.700 53.100 81.000 53.800 ;
        RECT 82.600 53.600 83.000 53.800 ;
        RECT 81.500 53.100 83.300 53.300 ;
        RECT 76.600 51.100 77.000 52.100 ;
        RECT 79.000 51.100 79.400 52.100 ;
        RECT 80.600 51.100 81.000 53.100 ;
        RECT 81.400 53.000 83.400 53.100 ;
        RECT 81.400 51.100 81.800 53.000 ;
        RECT 83.000 51.100 83.400 53.000 ;
        RECT 84.600 52.100 84.900 53.800 ;
        RECT 85.400 52.400 85.800 53.200 ;
        RECT 86.300 53.100 86.600 53.800 ;
        RECT 88.200 53.600 88.600 53.800 ;
        RECT 87.100 53.100 88.900 53.300 ;
        RECT 84.600 51.100 85.000 52.100 ;
        RECT 86.200 51.100 86.600 53.100 ;
        RECT 87.000 53.000 89.000 53.100 ;
        RECT 87.000 51.100 87.400 53.000 ;
        RECT 88.600 51.100 89.000 53.000 ;
        RECT 89.400 51.100 89.800 53.800 ;
        RECT 91.000 51.100 91.400 59.900 ;
        RECT 92.600 56.200 93.000 59.900 ;
        RECT 96.300 56.200 96.700 59.900 ;
        RECT 97.000 56.800 97.400 57.200 ;
        RECT 97.100 56.200 97.400 56.800 ;
        RECT 92.600 55.900 93.700 56.200 ;
        RECT 96.300 55.900 96.800 56.200 ;
        RECT 97.100 55.900 97.800 56.200 ;
        RECT 93.400 55.600 93.700 55.900 ;
        RECT 93.400 55.200 94.000 55.600 ;
        RECT 92.600 54.400 93.000 55.200 ;
        RECT 93.400 53.700 93.700 55.200 ;
        RECT 95.800 54.400 96.200 55.200 ;
        RECT 96.500 54.200 96.800 55.900 ;
        RECT 97.400 55.800 97.800 55.900 ;
        RECT 95.000 54.100 95.400 54.200 ;
        RECT 95.000 53.800 95.800 54.100 ;
        RECT 96.500 53.800 97.800 54.200 ;
        RECT 92.600 53.400 93.700 53.700 ;
        RECT 95.400 53.600 95.800 53.800 ;
        RECT 92.600 51.100 93.000 53.400 ;
        RECT 95.100 53.100 96.900 53.300 ;
        RECT 97.400 53.100 97.700 53.800 ;
        RECT 95.000 53.000 97.000 53.100 ;
        RECT 95.000 51.100 95.400 53.000 ;
        RECT 96.600 51.100 97.000 53.000 ;
        RECT 97.400 51.100 97.800 53.100 ;
        RECT 1.400 47.100 1.800 49.900 ;
        RECT 3.500 49.200 3.900 49.900 ;
        RECT 3.500 48.800 4.200 49.200 ;
        RECT 3.500 48.200 3.900 48.800 ;
        RECT 3.000 47.900 3.900 48.200 ;
        RECT 4.600 48.000 5.000 49.900 ;
        RECT 6.200 48.000 6.600 49.900 ;
        RECT 4.600 47.900 6.600 48.000 ;
        RECT 7.000 47.900 7.400 49.900 ;
        RECT 7.800 47.900 8.200 49.900 ;
        RECT 9.900 49.200 10.300 49.900 ;
        RECT 9.900 48.800 10.600 49.200 ;
        RECT 11.800 48.900 12.200 49.900 ;
        RECT 9.900 48.400 10.300 48.800 ;
        RECT 9.900 47.900 10.600 48.400 ;
        RECT 2.200 47.100 2.600 47.600 ;
        RECT 1.400 46.800 2.600 47.100 ;
        RECT 0.600 46.100 1.000 46.200 ;
        RECT 1.400 46.100 1.800 46.800 ;
        RECT 0.600 45.800 1.800 46.100 ;
        RECT 1.400 41.100 1.800 45.800 ;
        RECT 3.000 41.100 3.400 47.900 ;
        RECT 4.700 47.700 6.500 47.900 ;
        RECT 7.000 47.200 7.300 47.900 ;
        RECT 7.900 47.800 8.200 47.900 ;
        RECT 7.900 47.600 8.800 47.800 ;
        RECT 7.900 47.500 10.000 47.600 ;
        RECT 8.500 47.300 10.000 47.500 ;
        RECT 9.600 47.200 10.000 47.300 ;
        RECT 6.100 46.800 7.400 47.200 ;
        RECT 3.800 44.400 4.200 45.200 ;
        RECT 6.100 45.100 6.400 46.800 ;
        RECT 9.600 45.500 9.900 47.200 ;
        RECT 10.300 46.200 10.600 47.900 ;
        RECT 10.200 45.800 10.600 46.200 ;
        RECT 8.700 45.200 9.900 45.500 ;
        RECT 7.000 45.100 7.400 45.200 ;
        RECT 5.900 44.800 6.400 45.100 ;
        RECT 6.700 44.800 7.400 45.100 ;
        RECT 5.900 41.100 6.300 44.800 ;
        RECT 6.700 44.200 7.000 44.800 ;
        RECT 6.600 43.800 7.000 44.200 ;
        RECT 8.700 43.100 9.000 45.200 ;
        RECT 10.300 45.100 10.600 45.800 ;
        RECT 11.800 48.200 12.100 48.900 ;
        RECT 13.500 48.200 13.900 48.600 ;
        RECT 11.800 47.800 12.200 48.200 ;
        RECT 13.400 47.800 13.800 48.200 ;
        RECT 14.200 47.900 14.600 49.900 ;
        RECT 11.800 47.200 12.100 47.800 ;
        RECT 11.800 46.800 12.200 47.200 ;
        RECT 11.800 45.100 12.100 46.800 ;
        RECT 13.400 46.100 13.800 46.200 ;
        RECT 14.300 46.100 14.600 47.900 ;
        RECT 16.600 47.900 17.000 49.900 ;
        RECT 18.200 48.900 18.600 49.900 ;
        RECT 15.000 47.100 15.400 47.200 ;
        RECT 16.600 47.100 16.900 47.900 ;
        RECT 18.200 47.800 18.500 48.900 ;
        RECT 19.800 48.000 20.200 49.900 ;
        RECT 21.400 48.000 21.800 49.900 ;
        RECT 19.800 47.900 21.800 48.000 ;
        RECT 22.200 47.900 22.600 49.900 ;
        RECT 24.800 49.200 25.200 49.900 ;
        RECT 24.600 48.800 25.200 49.200 ;
        RECT 15.000 46.800 16.900 47.100 ;
        RECT 15.000 46.400 15.400 46.800 ;
        RECT 16.600 46.200 16.900 46.800 ;
        RECT 17.300 47.500 18.500 47.800 ;
        RECT 19.900 47.700 21.700 47.900 ;
        RECT 15.800 46.100 16.200 46.200 ;
        RECT 13.400 45.800 14.600 46.100 ;
        RECT 15.400 45.800 16.200 46.100 ;
        RECT 16.600 45.800 17.000 46.200 ;
        RECT 17.300 46.000 17.600 47.500 ;
        RECT 20.200 47.200 20.600 47.400 ;
        RECT 22.200 47.200 22.500 47.900 ;
        RECT 19.800 46.900 20.600 47.200 ;
        RECT 19.800 46.800 20.200 46.900 ;
        RECT 21.300 46.800 22.600 47.200 ;
        RECT 24.800 47.100 25.200 48.800 ;
        RECT 26.500 48.200 26.900 49.900 ;
        RECT 28.600 49.100 29.000 49.200 ;
        RECT 30.500 49.100 30.900 49.900 ;
        RECT 28.600 48.800 30.900 49.100 ;
        RECT 30.500 48.200 30.900 48.800 ;
        RECT 26.500 47.900 27.400 48.200 ;
        RECT 30.500 47.900 31.400 48.200 ;
        RECT 33.900 47.900 34.700 49.900 ;
        RECT 37.900 49.200 38.300 49.900 ;
        RECT 37.400 48.800 38.300 49.200 ;
        RECT 37.900 48.200 38.300 48.800 ;
        RECT 37.400 47.900 38.300 48.200 ;
        RECT 40.300 47.900 41.100 49.900 ;
        RECT 43.000 47.900 43.400 49.900 ;
        RECT 43.800 48.000 44.200 49.900 ;
        RECT 45.400 48.000 45.800 49.900 ;
        RECT 47.000 48.800 47.400 49.900 ;
        RECT 43.800 47.900 45.800 48.000 ;
        RECT 24.800 46.900 25.700 47.100 ;
        RECT 24.900 46.800 25.700 46.900 ;
        RECT 13.500 45.100 13.800 45.800 ;
        RECT 15.400 45.600 15.800 45.800 ;
        RECT 16.600 45.100 16.900 45.800 ;
        RECT 17.300 45.700 17.700 46.000 ;
        RECT 20.600 45.800 21.000 46.600 ;
        RECT 17.300 45.600 19.400 45.700 ;
        RECT 17.400 45.400 19.400 45.600 ;
        RECT 8.600 41.100 9.000 43.100 ;
        RECT 10.200 41.100 10.600 45.100 ;
        RECT 11.300 44.700 12.200 45.100 ;
        RECT 11.300 41.100 11.700 44.700 ;
        RECT 13.400 41.100 13.800 45.100 ;
        RECT 14.200 44.800 16.200 45.100 ;
        RECT 16.600 44.800 17.300 45.100 ;
        RECT 14.200 41.100 14.600 44.800 ;
        RECT 15.800 41.100 16.200 44.800 ;
        RECT 16.900 44.200 17.300 44.800 ;
        RECT 16.600 43.800 17.300 44.200 ;
        RECT 16.900 41.100 17.300 43.800 ;
        RECT 19.000 41.100 19.400 45.400 ;
        RECT 21.300 45.100 21.600 46.800 ;
        RECT 23.800 45.800 24.600 46.200 ;
        RECT 22.200 45.100 22.600 45.200 ;
        RECT 23.000 45.100 23.400 45.600 ;
        RECT 25.400 45.200 25.700 46.800 ;
        RECT 21.100 44.800 21.600 45.100 ;
        RECT 21.900 44.800 24.100 45.100 ;
        RECT 21.100 42.200 21.500 44.800 ;
        RECT 21.900 44.200 22.200 44.800 ;
        RECT 21.800 43.800 22.200 44.200 ;
        RECT 23.800 44.200 24.100 44.800 ;
        RECT 25.400 44.800 25.800 45.200 ;
        RECT 23.800 43.800 24.200 44.200 ;
        RECT 24.600 43.800 25.000 44.600 ;
        RECT 25.400 43.500 25.700 44.800 ;
        RECT 23.900 43.200 25.700 43.500 ;
        RECT 23.900 43.100 24.200 43.200 ;
        RECT 20.600 41.800 21.500 42.200 ;
        RECT 21.100 41.100 21.500 41.800 ;
        RECT 23.800 41.100 24.200 43.100 ;
        RECT 25.400 43.100 25.700 43.200 ;
        RECT 25.400 41.100 25.800 43.100 ;
        RECT 27.000 41.100 27.400 47.900 ;
        RECT 30.200 44.400 30.600 45.200 ;
        RECT 31.000 41.100 31.400 47.900 ;
        RECT 31.800 47.100 32.200 47.600 ;
        RECT 33.400 47.100 33.800 47.200 ;
        RECT 31.800 46.800 33.800 47.100 ;
        RECT 33.500 46.600 33.800 46.800 ;
        RECT 33.500 46.200 33.900 46.600 ;
        RECT 34.200 46.200 34.500 47.900 ;
        RECT 36.600 46.800 37.000 47.600 ;
        RECT 32.600 45.400 33.000 46.200 ;
        RECT 34.200 45.800 34.600 46.200 ;
        RECT 35.800 46.100 36.200 46.200 ;
        RECT 35.400 45.800 36.200 46.100 ;
        RECT 34.200 45.700 34.500 45.800 ;
        RECT 33.500 45.400 34.500 45.700 ;
        RECT 35.400 45.600 35.800 45.800 ;
        RECT 33.500 45.100 33.800 45.400 ;
        RECT 32.600 41.400 33.000 45.100 ;
        RECT 33.400 41.700 33.800 45.100 ;
        RECT 34.200 44.800 36.200 45.100 ;
        RECT 34.200 41.400 34.600 44.800 ;
        RECT 32.600 41.100 34.600 41.400 ;
        RECT 35.800 41.100 36.200 44.800 ;
        RECT 37.400 41.100 37.800 47.900 ;
        RECT 39.800 46.800 40.200 47.200 ;
        RECT 39.900 46.600 40.200 46.800 ;
        RECT 39.900 46.200 40.300 46.600 ;
        RECT 40.600 46.200 40.900 47.900 ;
        RECT 43.100 47.200 43.400 47.900 ;
        RECT 43.900 47.700 45.700 47.900 ;
        RECT 46.200 47.800 46.600 48.600 ;
        RECT 45.000 47.200 45.400 47.400 ;
        RECT 47.100 47.200 47.400 48.800 ;
        RECT 43.000 46.800 44.300 47.200 ;
        RECT 45.000 46.900 45.800 47.200 ;
        RECT 45.400 46.800 45.800 46.900 ;
        RECT 47.000 46.800 47.400 47.200 ;
        RECT 48.600 46.800 49.000 47.600 ;
        RECT 39.000 45.400 39.400 46.200 ;
        RECT 40.600 45.800 41.000 46.200 ;
        RECT 42.200 46.100 42.600 46.200 ;
        RECT 41.800 45.800 42.600 46.100 ;
        RECT 40.600 45.700 40.900 45.800 ;
        RECT 39.900 45.400 40.900 45.700 ;
        RECT 41.800 45.600 42.200 45.800 ;
        RECT 38.200 44.400 38.600 45.200 ;
        RECT 39.900 45.100 40.200 45.400 ;
        RECT 43.000 45.100 43.400 45.200 ;
        RECT 44.000 45.100 44.300 46.800 ;
        RECT 44.600 45.800 45.000 46.600 ;
        RECT 47.100 45.100 47.400 46.800 ;
        RECT 47.800 45.400 48.200 46.200 ;
        RECT 39.000 41.400 39.400 45.100 ;
        RECT 39.800 41.700 40.200 45.100 ;
        RECT 40.600 44.800 42.600 45.100 ;
        RECT 43.000 44.800 43.700 45.100 ;
        RECT 44.000 44.800 44.500 45.100 ;
        RECT 40.600 41.400 41.000 44.800 ;
        RECT 39.000 41.100 41.000 41.400 ;
        RECT 42.200 41.100 42.600 44.800 ;
        RECT 43.400 44.200 43.700 44.800 ;
        RECT 43.400 43.800 43.800 44.200 ;
        RECT 44.100 41.100 44.500 44.800 ;
        RECT 47.000 44.700 47.900 45.100 ;
        RECT 47.500 41.100 47.900 44.700 ;
        RECT 49.400 41.100 49.800 49.900 ;
        RECT 50.200 41.100 50.600 49.900 ;
        RECT 51.800 47.900 52.200 49.900 ;
        RECT 52.600 48.000 53.000 49.900 ;
        RECT 54.200 48.000 54.600 49.900 ;
        RECT 55.100 48.200 55.500 48.600 ;
        RECT 52.600 47.900 54.600 48.000 ;
        RECT 51.000 46.800 51.400 47.600 ;
        RECT 51.900 47.200 52.200 47.900 ;
        RECT 52.700 47.700 54.500 47.900 ;
        RECT 55.000 47.800 55.400 48.200 ;
        RECT 55.800 47.900 56.200 49.900 ;
        RECT 53.800 47.200 54.200 47.400 ;
        RECT 51.800 46.800 53.100 47.200 ;
        RECT 53.800 46.900 54.600 47.200 ;
        RECT 54.200 46.800 54.600 46.900 ;
        RECT 51.800 45.100 52.200 45.200 ;
        RECT 52.800 45.100 53.100 46.800 ;
        RECT 53.400 45.800 53.800 46.600 ;
        RECT 55.000 46.100 55.400 46.200 ;
        RECT 55.900 46.100 56.200 47.900 ;
        RECT 56.600 46.400 57.000 47.200 ;
        RECT 60.000 47.100 60.400 49.900 ;
        RECT 61.400 48.000 61.800 49.900 ;
        RECT 63.000 48.000 63.400 49.900 ;
        RECT 61.400 47.900 63.400 48.000 ;
        RECT 63.800 47.900 64.200 49.900 ;
        RECT 64.600 48.000 65.000 49.900 ;
        RECT 66.200 48.000 66.600 49.900 ;
        RECT 64.600 47.900 66.600 48.000 ;
        RECT 67.000 47.900 67.400 49.900 ;
        RECT 71.000 47.900 71.400 49.900 ;
        RECT 71.700 48.200 72.100 48.600 ;
        RECT 61.500 47.700 63.300 47.900 ;
        RECT 61.800 47.200 62.200 47.400 ;
        RECT 63.800 47.200 64.100 47.900 ;
        RECT 64.700 47.700 66.500 47.900 ;
        RECT 65.000 47.200 65.400 47.400 ;
        RECT 67.000 47.200 67.300 47.900 ;
        RECT 60.000 46.900 60.900 47.100 ;
        RECT 60.100 46.800 60.900 46.900 ;
        RECT 61.400 46.900 62.200 47.200 ;
        RECT 61.400 46.800 61.800 46.900 ;
        RECT 62.900 46.800 64.200 47.200 ;
        RECT 64.600 46.900 65.400 47.200 ;
        RECT 64.600 46.800 65.000 46.900 ;
        RECT 66.100 46.800 67.400 47.200 ;
        RECT 60.600 46.200 60.900 46.800 ;
        RECT 55.000 45.800 56.200 46.100 ;
        RECT 59.000 45.800 59.800 46.200 ;
        RECT 60.600 45.800 61.000 46.200 ;
        RECT 62.200 45.800 62.600 46.600 ;
        RECT 55.100 45.100 55.400 45.800 ;
        RECT 58.200 45.100 58.600 45.600 ;
        RECT 60.600 45.200 60.900 45.800 ;
        RECT 59.000 45.100 59.400 45.200 ;
        RECT 51.800 44.800 52.500 45.100 ;
        RECT 52.800 44.800 53.300 45.100 ;
        RECT 52.200 44.200 52.500 44.800 ;
        RECT 52.200 43.800 52.600 44.200 ;
        RECT 52.900 41.100 53.300 44.800 ;
        RECT 55.000 41.100 55.400 45.100 ;
        RECT 55.800 44.800 57.800 45.100 ;
        RECT 58.200 44.800 59.400 45.100 ;
        RECT 60.600 44.800 61.000 45.200 ;
        RECT 62.900 45.100 63.200 46.800 ;
        RECT 63.800 45.800 64.200 46.200 ;
        RECT 65.400 45.800 65.800 46.600 ;
        RECT 66.100 46.100 66.400 46.800 ;
        RECT 70.200 46.400 70.600 47.200 ;
        RECT 67.800 46.100 68.200 46.200 ;
        RECT 66.100 45.800 68.200 46.100 ;
        RECT 69.400 46.100 69.800 46.200 ;
        RECT 71.000 46.100 71.300 47.900 ;
        RECT 71.800 47.800 72.200 48.200 ;
        RECT 74.400 47.100 74.800 49.900 ;
        RECT 74.400 46.900 75.300 47.100 ;
        RECT 74.500 46.800 75.300 46.900 ;
        RECT 75.800 46.800 76.200 47.600 ;
        RECT 71.800 46.100 72.200 46.200 ;
        RECT 69.400 45.800 70.200 46.100 ;
        RECT 71.000 45.800 72.200 46.100 ;
        RECT 73.400 45.800 74.200 46.200 ;
        RECT 63.800 45.200 64.100 45.800 ;
        RECT 63.800 45.100 64.200 45.200 ;
        RECT 66.100 45.100 66.400 45.800 ;
        RECT 69.800 45.600 70.200 45.800 ;
        RECT 67.000 45.100 67.400 45.200 ;
        RECT 71.800 45.100 72.100 45.800 ;
        RECT 62.700 44.800 63.200 45.100 ;
        RECT 63.500 44.800 64.200 45.100 ;
        RECT 65.900 44.800 66.400 45.100 ;
        RECT 66.700 44.800 67.400 45.100 ;
        RECT 69.400 44.800 71.400 45.100 ;
        RECT 55.800 41.100 56.200 44.800 ;
        RECT 57.400 41.100 57.800 44.800 ;
        RECT 59.800 43.800 60.200 44.600 ;
        RECT 60.600 43.500 60.900 44.800 ;
        RECT 59.100 43.200 60.900 43.500 ;
        RECT 59.100 43.100 59.400 43.200 ;
        RECT 59.000 41.100 59.400 43.100 ;
        RECT 60.600 43.100 60.900 43.200 ;
        RECT 60.600 41.100 61.000 43.100 ;
        RECT 62.700 41.100 63.100 44.800 ;
        RECT 63.500 44.200 63.800 44.800 ;
        RECT 63.400 43.800 63.800 44.200 ;
        RECT 65.900 41.100 66.300 44.800 ;
        RECT 66.700 44.200 67.000 44.800 ;
        RECT 66.600 43.800 67.000 44.200 ;
        RECT 69.400 41.100 69.800 44.800 ;
        RECT 71.000 41.100 71.400 44.800 ;
        RECT 71.800 41.100 72.200 45.100 ;
        RECT 72.600 44.800 73.000 45.600 ;
        RECT 75.000 45.200 75.300 46.800 ;
        RECT 75.000 44.800 75.400 45.200 ;
        RECT 74.200 43.800 74.600 44.600 ;
        RECT 75.000 43.500 75.300 44.800 ;
        RECT 73.500 43.200 75.300 43.500 ;
        RECT 73.500 43.100 73.800 43.200 ;
        RECT 73.400 41.100 73.800 43.100 ;
        RECT 75.000 41.100 75.400 43.200 ;
        RECT 76.600 41.100 77.000 49.900 ;
        RECT 77.400 48.000 77.800 49.900 ;
        RECT 79.000 48.000 79.400 49.900 ;
        RECT 77.400 47.900 79.400 48.000 ;
        RECT 79.800 47.900 80.200 49.900 ;
        RECT 82.200 47.900 82.600 49.900 ;
        RECT 84.600 48.900 85.000 49.900 ;
        RECT 88.600 48.900 89.000 49.900 ;
        RECT 90.200 49.200 90.600 49.900 ;
        RECT 82.900 48.200 83.300 48.600 ;
        RECT 77.500 47.700 79.300 47.900 ;
        RECT 77.800 47.200 78.200 47.400 ;
        RECT 79.800 47.200 80.100 47.900 ;
        RECT 77.400 46.900 78.200 47.200 ;
        RECT 77.400 46.800 77.800 46.900 ;
        RECT 78.900 46.800 80.200 47.200 ;
        RECT 78.200 45.800 78.600 46.600 ;
        RECT 78.900 46.200 79.200 46.800 ;
        RECT 81.400 46.400 81.800 47.200 ;
        RECT 78.900 45.800 79.400 46.200 ;
        RECT 80.600 46.100 81.000 46.200 ;
        RECT 82.200 46.100 82.500 47.900 ;
        RECT 83.000 47.800 83.400 48.200 ;
        RECT 83.800 47.800 84.200 48.600 ;
        RECT 83.000 47.100 83.300 47.800 ;
        RECT 84.700 47.200 85.000 48.900 ;
        RECT 88.400 48.800 89.000 48.900 ;
        RECT 90.100 48.800 90.600 49.200 ;
        RECT 88.400 48.500 90.400 48.800 ;
        RECT 83.800 47.100 84.200 47.200 ;
        RECT 83.000 46.800 84.200 47.100 ;
        RECT 84.600 47.100 85.000 47.200 ;
        RECT 85.400 47.100 85.800 47.200 ;
        RECT 84.600 46.800 85.800 47.100 ;
        RECT 83.000 46.100 83.400 46.200 ;
        RECT 80.600 45.800 81.400 46.100 ;
        RECT 82.200 45.800 83.400 46.100 ;
        RECT 78.900 45.100 79.200 45.800 ;
        RECT 81.000 45.600 81.400 45.800 ;
        RECT 79.800 45.100 80.200 45.200 ;
        RECT 83.000 45.100 83.300 45.800 ;
        RECT 84.700 45.100 85.000 46.800 ;
        RECT 85.400 45.400 85.800 46.200 ;
        RECT 88.400 45.200 88.700 48.500 ;
        RECT 90.200 47.800 91.400 48.200 ;
        RECT 92.600 47.600 93.000 49.900 ;
        RECT 95.000 47.900 95.400 49.900 ;
        RECT 97.100 49.200 97.500 49.900 ;
        RECT 97.100 48.800 97.800 49.200 ;
        RECT 97.100 48.400 97.500 48.800 ;
        RECT 97.100 47.900 97.800 48.400 ;
        RECT 95.100 47.800 95.400 47.900 ;
        RECT 95.100 47.600 96.000 47.800 ;
        RECT 92.600 47.300 93.700 47.600 ;
        RECT 95.100 47.500 97.200 47.600 ;
        RECT 95.700 47.300 97.200 47.500 ;
        RECT 89.800 47.100 90.600 47.200 ;
        RECT 91.000 47.100 91.400 47.200 ;
        RECT 89.800 46.800 91.400 47.100 ;
        RECT 89.000 45.800 89.800 46.200 ;
        RECT 90.200 46.100 90.600 46.200 ;
        RECT 92.600 46.100 93.000 46.600 ;
        RECT 90.200 45.800 93.000 46.100 ;
        RECT 93.400 45.800 93.700 47.300 ;
        RECT 96.800 47.200 97.200 47.300 ;
        RECT 95.000 45.800 95.400 47.200 ;
        RECT 96.000 46.900 96.400 47.000 ;
        RECT 95.900 46.600 96.400 46.900 ;
        RECT 95.900 46.200 96.200 46.600 ;
        RECT 95.800 45.800 96.200 46.200 ;
        RECT 78.700 44.800 79.200 45.100 ;
        RECT 79.500 44.800 80.200 45.100 ;
        RECT 80.600 44.800 82.600 45.100 ;
        RECT 78.700 41.100 79.100 44.800 ;
        RECT 79.500 44.200 79.800 44.800 ;
        RECT 79.400 43.800 79.800 44.200 ;
        RECT 80.600 41.100 81.000 44.800 ;
        RECT 82.200 41.100 82.600 44.800 ;
        RECT 83.000 41.100 83.400 45.100 ;
        RECT 84.600 44.700 85.500 45.100 ;
        RECT 87.000 44.900 88.700 45.200 ;
        RECT 93.400 45.400 94.000 45.800 ;
        RECT 96.800 45.500 97.100 47.200 ;
        RECT 97.500 46.200 97.800 47.900 ;
        RECT 97.400 45.800 97.800 46.200 ;
        RECT 93.400 45.100 93.700 45.400 ;
        RECT 87.000 44.800 87.400 44.900 ;
        RECT 85.100 41.100 85.500 44.700 ;
        RECT 87.100 44.500 87.400 44.800 ;
        RECT 92.600 44.800 93.700 45.100 ;
        RECT 95.900 45.200 97.100 45.500 ;
        RECT 87.900 44.500 89.700 44.600 ;
        RECT 86.200 41.500 86.600 44.500 ;
        RECT 87.000 41.700 87.400 44.500 ;
        RECT 87.800 44.300 89.700 44.500 ;
        RECT 86.300 41.400 86.600 41.500 ;
        RECT 87.800 41.500 88.200 44.300 ;
        RECT 89.400 44.100 89.700 44.300 ;
        RECT 90.300 44.400 92.100 44.700 ;
        RECT 90.300 44.100 90.600 44.400 ;
        RECT 87.800 41.400 88.100 41.500 ;
        RECT 86.300 41.100 88.100 41.400 ;
        RECT 88.600 41.400 89.000 44.000 ;
        RECT 89.400 41.700 89.800 44.100 ;
        RECT 90.200 41.400 90.600 44.100 ;
        RECT 88.600 41.100 90.600 41.400 ;
        RECT 91.800 44.100 92.100 44.400 ;
        RECT 91.800 41.100 92.200 44.100 ;
        RECT 92.600 41.100 93.000 44.800 ;
        RECT 95.900 43.100 96.200 45.200 ;
        RECT 97.500 45.100 97.800 45.800 ;
        RECT 95.800 41.100 96.200 43.100 ;
        RECT 97.400 41.100 97.800 45.100 ;
        RECT 1.900 36.200 2.300 39.900 ;
        RECT 2.600 36.800 3.000 37.200 ;
        RECT 2.700 36.200 3.000 36.800 ;
        RECT 3.800 36.200 4.200 39.900 ;
        RECT 5.400 39.600 7.400 39.900 ;
        RECT 5.400 36.200 5.800 39.600 ;
        RECT 1.900 35.900 2.400 36.200 ;
        RECT 2.700 35.900 3.400 36.200 ;
        RECT 3.800 35.900 5.800 36.200 ;
        RECT 6.200 35.900 6.600 39.300 ;
        RECT 7.000 35.900 7.400 39.600 ;
        RECT 1.400 34.400 1.800 35.200 ;
        RECT 2.100 34.200 2.400 35.900 ;
        RECT 3.000 35.800 3.400 35.900 ;
        RECT 6.200 35.600 6.500 35.900 ;
        RECT 4.200 35.200 4.600 35.400 ;
        RECT 5.500 35.300 6.500 35.600 ;
        RECT 5.500 35.200 5.800 35.300 ;
        RECT 3.800 34.900 4.600 35.200 ;
        RECT 3.800 34.800 4.200 34.900 ;
        RECT 5.400 34.800 5.800 35.200 ;
        RECT 7.000 34.800 7.400 35.600 ;
        RECT 3.800 34.200 4.100 34.800 ;
        RECT 0.600 34.100 1.000 34.200 ;
        RECT 0.600 33.800 1.400 34.100 ;
        RECT 2.100 33.800 3.400 34.200 ;
        RECT 3.800 33.800 4.200 34.200 ;
        RECT 4.600 33.800 5.000 34.600 ;
        RECT 1.000 33.600 1.400 33.800 ;
        RECT 0.700 33.100 2.500 33.300 ;
        RECT 3.000 33.100 3.300 33.800 ;
        RECT 5.500 33.100 5.800 34.800 ;
        RECT 6.100 34.400 6.500 34.800 ;
        RECT 6.200 34.200 6.500 34.400 ;
        RECT 6.200 33.800 6.600 34.200 ;
        RECT 0.600 33.000 2.600 33.100 ;
        RECT 0.600 31.100 1.000 33.000 ;
        RECT 2.200 31.100 2.600 33.000 ;
        RECT 3.000 31.100 3.400 33.100 ;
        RECT 5.300 31.100 6.100 33.100 ;
        RECT 8.600 31.100 9.000 39.900 ;
        RECT 10.700 36.200 11.100 39.900 ;
        RECT 11.400 36.800 11.800 37.200 ;
        RECT 11.500 36.200 11.800 36.800 ;
        RECT 13.900 36.300 14.300 39.900 ;
        RECT 10.700 35.900 11.200 36.200 ;
        RECT 11.500 35.900 12.200 36.200 ;
        RECT 13.400 35.900 14.300 36.300 ;
        RECT 10.900 34.200 11.200 35.900 ;
        RECT 11.800 35.800 12.200 35.900 ;
        RECT 13.500 34.200 13.800 35.900 ;
        RECT 15.000 35.600 15.400 39.900 ;
        RECT 17.100 36.200 17.500 39.900 ;
        RECT 18.200 36.200 18.600 39.900 ;
        RECT 19.800 36.200 20.200 39.900 ;
        RECT 17.100 35.900 17.800 36.200 ;
        RECT 18.200 35.900 20.200 36.200 ;
        RECT 20.600 35.900 21.000 39.900 ;
        RECT 21.400 36.200 21.800 39.900 ;
        RECT 23.000 36.200 23.400 39.900 ;
        RECT 21.400 35.900 23.400 36.200 ;
        RECT 23.800 35.900 24.200 39.900 ;
        RECT 24.900 36.300 25.300 39.900 ;
        RECT 24.900 35.900 25.800 36.300 ;
        RECT 29.900 36.200 30.300 39.900 ;
        RECT 30.600 36.800 31.000 37.200 ;
        RECT 30.700 36.200 31.000 36.800 ;
        RECT 29.900 35.900 30.400 36.200 ;
        RECT 30.700 35.900 31.400 36.200 ;
        RECT 14.200 34.800 14.600 35.600 ;
        RECT 15.000 35.400 17.000 35.600 ;
        RECT 15.000 35.300 17.100 35.400 ;
        RECT 16.700 35.000 17.100 35.300 ;
        RECT 17.500 35.200 17.800 35.900 ;
        RECT 18.600 35.200 19.000 35.400 ;
        RECT 20.600 35.200 20.900 35.900 ;
        RECT 21.800 35.200 22.200 35.400 ;
        RECT 23.800 35.200 24.100 35.900 ;
        RECT 9.400 34.100 9.800 34.200 ;
        RECT 9.400 33.800 10.200 34.100 ;
        RECT 10.900 33.800 12.200 34.200 ;
        RECT 13.400 33.800 13.800 34.200 ;
        RECT 9.800 33.600 10.200 33.800 ;
        RECT 9.500 33.100 11.300 33.300 ;
        RECT 11.800 33.100 12.100 33.800 ;
        RECT 9.400 33.000 11.400 33.100 ;
        RECT 9.400 31.100 9.800 33.000 ;
        RECT 11.000 31.100 11.400 33.000 ;
        RECT 11.800 31.100 12.200 33.100 ;
        RECT 13.500 32.200 13.800 33.800 ;
        RECT 16.800 33.500 17.100 35.000 ;
        RECT 17.400 35.100 17.800 35.200 ;
        RECT 18.200 35.100 19.000 35.200 ;
        RECT 17.400 34.900 19.000 35.100 ;
        RECT 19.800 34.900 21.000 35.200 ;
        RECT 17.400 34.800 18.600 34.900 ;
        RECT 15.900 33.200 17.100 33.500 ;
        RECT 15.000 32.400 15.400 33.200 ;
        RECT 13.400 31.100 13.800 32.200 ;
        RECT 15.900 32.100 16.200 33.200 ;
        RECT 17.500 33.100 17.800 34.800 ;
        RECT 18.200 34.200 18.500 34.800 ;
        RECT 18.200 33.800 18.600 34.200 ;
        RECT 19.000 33.800 19.400 34.600 ;
        RECT 15.800 31.100 16.200 32.100 ;
        RECT 17.400 31.100 17.800 33.100 ;
        RECT 19.800 33.100 20.100 34.900 ;
        RECT 20.600 34.800 21.000 34.900 ;
        RECT 21.400 34.900 22.200 35.200 ;
        RECT 23.000 34.900 24.200 35.200 ;
        RECT 21.400 34.800 21.800 34.900 ;
        RECT 22.200 33.800 22.600 34.600 ;
        RECT 23.000 34.100 23.300 34.900 ;
        RECT 23.800 34.800 24.200 34.900 ;
        RECT 24.600 34.800 25.000 35.600 ;
        RECT 25.400 35.100 25.700 35.900 ;
        RECT 29.400 35.100 29.800 35.200 ;
        RECT 25.400 34.800 29.800 35.100 ;
        RECT 25.400 34.200 25.700 34.800 ;
        RECT 29.400 34.400 29.800 34.800 ;
        RECT 30.100 35.100 30.400 35.900 ;
        RECT 31.000 35.800 31.400 35.900 ;
        RECT 31.800 35.800 32.200 36.600 ;
        RECT 31.800 35.100 32.100 35.800 ;
        RECT 30.100 34.800 32.100 35.100 ;
        RECT 30.100 34.200 30.400 34.800 ;
        RECT 23.800 34.100 24.200 34.200 ;
        RECT 23.000 33.800 24.200 34.100 ;
        RECT 25.400 33.800 25.800 34.200 ;
        RECT 27.000 34.100 27.400 34.200 ;
        RECT 28.600 34.100 29.000 34.200 ;
        RECT 27.000 33.800 29.400 34.100 ;
        RECT 30.100 33.800 31.400 34.200 ;
        RECT 19.800 31.100 20.200 33.100 ;
        RECT 20.600 32.800 21.000 33.200 ;
        RECT 23.000 33.100 23.300 33.800 ;
        RECT 20.500 32.400 20.900 32.800 ;
        RECT 23.000 31.100 23.400 33.100 ;
        RECT 23.800 32.800 24.200 33.200 ;
        RECT 23.700 32.400 24.100 32.800 ;
        RECT 25.400 32.100 25.700 33.800 ;
        RECT 29.000 33.600 29.400 33.800 ;
        RECT 28.700 33.100 30.500 33.300 ;
        RECT 31.000 33.100 31.300 33.800 ;
        RECT 32.600 33.100 33.000 39.900 ;
        RECT 34.200 36.200 34.600 39.900 ;
        RECT 35.800 36.200 36.200 39.900 ;
        RECT 34.200 35.900 36.200 36.200 ;
        RECT 36.600 35.900 37.000 39.900 ;
        RECT 38.700 39.200 39.100 39.900 ;
        RECT 38.200 38.800 39.100 39.200 ;
        RECT 38.700 36.200 39.100 38.800 ;
        RECT 39.400 36.800 39.800 37.200 ;
        RECT 39.500 36.200 39.800 36.800 ;
        RECT 38.700 35.900 39.200 36.200 ;
        RECT 39.500 36.100 40.200 36.200 ;
        RECT 40.600 36.100 41.000 39.900 ;
        RECT 43.500 39.200 43.900 39.900 ;
        RECT 45.900 39.200 46.300 39.900 ;
        RECT 43.500 38.800 44.200 39.200 ;
        RECT 45.400 38.800 46.300 39.200 ;
        RECT 43.500 36.300 43.900 38.800 ;
        RECT 39.500 35.900 41.000 36.100 ;
        RECT 43.000 35.900 43.900 36.300 ;
        RECT 45.900 36.200 46.300 38.800 ;
        RECT 46.600 36.800 47.400 37.200 ;
        RECT 46.700 36.200 47.000 36.800 ;
        RECT 48.100 36.300 48.500 39.900 ;
        RECT 45.900 35.900 46.400 36.200 ;
        RECT 46.700 35.900 47.400 36.200 ;
        RECT 48.100 35.900 49.000 36.300 ;
        RECT 50.200 36.200 50.600 39.900 ;
        RECT 51.800 39.600 53.800 39.900 ;
        RECT 51.800 36.200 52.200 39.600 ;
        RECT 50.200 35.900 52.200 36.200 ;
        RECT 52.600 35.900 53.000 39.300 ;
        RECT 53.400 35.900 53.800 39.600 ;
        RECT 54.600 36.800 55.000 37.200 ;
        RECT 54.600 36.200 54.900 36.800 ;
        RECT 55.300 36.200 55.700 39.900 ;
        RECT 54.200 35.900 54.900 36.200 ;
        RECT 55.200 35.900 55.700 36.200 ;
        RECT 34.600 35.200 35.000 35.400 ;
        RECT 36.600 35.200 36.900 35.900 ;
        RECT 34.200 34.900 35.000 35.200 ;
        RECT 35.800 34.900 37.000 35.200 ;
        RECT 34.200 34.800 34.600 34.900 ;
        RECT 33.400 33.400 33.800 34.200 ;
        RECT 35.000 33.800 35.400 34.600 ;
        RECT 28.600 33.000 30.600 33.100 ;
        RECT 25.400 31.100 25.800 32.100 ;
        RECT 28.600 31.100 29.000 33.000 ;
        RECT 30.200 31.100 30.600 33.000 ;
        RECT 31.000 31.100 31.400 33.100 ;
        RECT 32.100 32.800 33.000 33.100 ;
        RECT 35.800 33.100 36.100 34.900 ;
        RECT 36.600 34.800 37.000 34.900 ;
        RECT 38.200 34.400 38.600 35.200 ;
        RECT 38.900 34.200 39.200 35.900 ;
        RECT 39.800 35.800 41.000 35.900 ;
        RECT 37.400 34.100 37.800 34.200 ;
        RECT 37.400 33.800 38.200 34.100 ;
        RECT 38.900 33.800 40.200 34.200 ;
        RECT 37.800 33.600 38.200 33.800 ;
        RECT 32.100 32.200 32.500 32.800 ;
        RECT 32.100 31.800 33.000 32.200 ;
        RECT 32.100 31.100 32.500 31.800 ;
        RECT 35.800 31.100 36.200 33.100 ;
        RECT 36.600 32.800 37.000 33.200 ;
        RECT 37.500 33.100 39.300 33.300 ;
        RECT 39.800 33.100 40.100 33.800 ;
        RECT 37.400 33.000 39.400 33.100 ;
        RECT 36.500 32.400 36.900 32.800 ;
        RECT 37.400 31.100 37.800 33.000 ;
        RECT 39.000 31.100 39.400 33.000 ;
        RECT 39.800 31.100 40.200 33.100 ;
        RECT 40.600 31.100 41.000 35.800 ;
        RECT 43.100 34.200 43.400 35.900 ;
        RECT 43.000 33.800 43.400 34.200 ;
        RECT 41.400 32.400 41.800 33.200 ;
        RECT 42.200 32.400 42.600 33.200 ;
        RECT 43.100 32.100 43.400 33.800 ;
        RECT 43.800 34.800 44.200 35.600 ;
        RECT 44.600 35.100 45.000 35.200 ;
        RECT 45.400 35.100 45.800 35.200 ;
        RECT 44.600 34.800 45.800 35.100 ;
        RECT 43.800 34.100 44.100 34.800 ;
        RECT 45.400 34.400 45.800 34.800 ;
        RECT 46.100 34.200 46.400 35.900 ;
        RECT 47.000 35.800 47.400 35.900 ;
        RECT 47.800 34.800 48.200 35.600 ;
        RECT 48.600 34.200 48.900 35.900 ;
        RECT 52.600 35.600 52.900 35.900 ;
        RECT 54.200 35.800 54.600 35.900 ;
        RECT 50.600 35.200 51.000 35.400 ;
        RECT 51.900 35.300 52.900 35.600 ;
        RECT 51.900 35.200 52.200 35.300 ;
        RECT 50.200 34.900 51.000 35.200 ;
        RECT 50.200 34.800 50.600 34.900 ;
        RECT 51.800 34.800 52.200 35.200 ;
        RECT 53.400 34.800 53.800 35.600 ;
        RECT 44.600 34.100 45.000 34.200 ;
        RECT 43.800 33.800 45.400 34.100 ;
        RECT 46.100 33.800 47.400 34.200 ;
        RECT 48.600 33.800 49.000 34.200 ;
        RECT 43.800 33.200 44.100 33.800 ;
        RECT 45.000 33.600 45.400 33.800 ;
        RECT 43.800 32.800 44.200 33.200 ;
        RECT 44.700 33.100 46.500 33.300 ;
        RECT 47.000 33.100 47.300 33.800 ;
        RECT 48.600 33.200 48.900 33.800 ;
        RECT 44.600 33.000 46.600 33.100 ;
        RECT 43.000 31.100 43.400 32.100 ;
        RECT 44.600 31.100 45.000 33.000 ;
        RECT 46.200 31.100 46.600 33.000 ;
        RECT 47.000 31.100 47.400 33.100 ;
        RECT 48.600 32.800 49.000 33.200 ;
        RECT 48.600 32.100 48.900 32.800 ;
        RECT 49.400 32.400 49.800 33.200 ;
        RECT 51.900 33.100 52.200 34.800 ;
        RECT 52.500 34.400 52.900 34.800 ;
        RECT 52.600 34.200 52.900 34.400 ;
        RECT 55.200 34.200 55.500 35.900 ;
        RECT 55.800 34.400 56.200 35.200 ;
        RECT 56.600 35.100 57.000 35.200 ;
        RECT 57.400 35.100 57.800 39.900 ;
        RECT 59.100 39.600 60.900 39.900 ;
        RECT 59.100 39.500 59.400 39.600 ;
        RECT 59.000 36.500 59.400 39.500 ;
        RECT 60.600 39.500 60.900 39.600 ;
        RECT 61.400 39.600 63.400 39.900 ;
        RECT 59.800 36.500 60.200 39.300 ;
        RECT 60.600 36.700 61.000 39.500 ;
        RECT 61.400 37.000 61.800 39.600 ;
        RECT 62.200 36.900 62.600 39.300 ;
        RECT 63.000 36.900 63.400 39.600 ;
        RECT 62.200 36.700 62.500 36.900 ;
        RECT 60.600 36.500 62.500 36.700 ;
        RECT 59.900 36.200 60.200 36.500 ;
        RECT 60.700 36.400 62.500 36.500 ;
        RECT 63.100 36.600 63.400 36.900 ;
        RECT 64.600 36.900 65.000 39.900 ;
        RECT 64.600 36.600 64.900 36.900 ;
        RECT 63.100 36.300 64.900 36.600 ;
        RECT 59.800 36.100 60.200 36.200 ;
        RECT 66.700 36.200 67.100 39.900 ;
        RECT 67.400 36.800 67.800 37.200 ;
        RECT 67.500 36.200 67.800 36.800 ;
        RECT 70.600 36.800 71.000 37.200 ;
        RECT 70.600 36.200 70.900 36.800 ;
        RECT 71.300 36.200 71.700 39.900 ;
        RECT 59.800 35.800 61.500 36.100 ;
        RECT 66.700 35.900 67.200 36.200 ;
        RECT 67.500 35.900 68.200 36.200 ;
        RECT 56.600 34.800 57.800 35.100 ;
        RECT 52.600 33.800 53.000 34.200 ;
        RECT 54.200 33.800 55.500 34.200 ;
        RECT 56.600 34.100 57.000 34.200 ;
        RECT 56.200 33.800 57.000 34.100 ;
        RECT 54.300 33.100 54.600 33.800 ;
        RECT 56.200 33.600 56.600 33.800 ;
        RECT 55.100 33.100 56.900 33.300 ;
        RECT 48.600 31.100 49.000 32.100 ;
        RECT 51.700 31.100 52.500 33.100 ;
        RECT 54.200 31.100 54.600 33.100 ;
        RECT 55.000 33.000 57.000 33.100 ;
        RECT 55.000 31.100 55.400 33.000 ;
        RECT 56.600 31.100 57.000 33.000 ;
        RECT 57.400 31.100 57.800 34.800 ;
        RECT 61.200 32.500 61.500 35.800 ;
        RECT 61.800 34.800 62.600 35.200 ;
        RECT 66.200 34.400 66.600 35.200 ;
        RECT 66.900 34.200 67.200 35.900 ;
        RECT 67.800 35.800 68.200 35.900 ;
        RECT 70.200 35.900 70.900 36.200 ;
        RECT 71.200 35.900 71.700 36.200 ;
        RECT 70.200 35.800 70.600 35.900 ;
        RECT 67.800 35.100 68.100 35.800 ;
        RECT 71.200 35.100 71.500 35.900 ;
        RECT 67.800 34.800 71.500 35.100 ;
        RECT 71.200 34.200 71.500 34.800 ;
        RECT 62.600 33.800 63.400 34.200 ;
        RECT 63.800 34.100 64.200 34.200 ;
        RECT 65.400 34.100 65.800 34.200 ;
        RECT 63.800 33.800 66.200 34.100 ;
        RECT 66.900 33.800 68.200 34.200 ;
        RECT 70.200 33.800 71.500 34.200 ;
        RECT 65.800 33.600 66.200 33.800 ;
        RECT 63.300 32.800 64.200 33.200 ;
        RECT 65.500 33.100 67.300 33.300 ;
        RECT 67.800 33.100 68.100 33.800 ;
        RECT 70.300 33.100 70.600 33.800 ;
        RECT 71.100 33.100 72.900 33.300 ;
        RECT 74.200 33.100 74.600 39.900 ;
        RECT 77.100 39.200 77.500 39.900 ;
        RECT 76.600 38.800 77.500 39.200 ;
        RECT 77.100 36.200 77.500 38.800 ;
        RECT 77.800 36.800 78.200 37.200 ;
        RECT 77.900 36.200 78.200 36.800 ;
        RECT 77.100 35.900 77.600 36.200 ;
        RECT 77.900 35.900 78.600 36.200 ;
        RECT 76.600 34.400 77.000 35.200 ;
        RECT 77.300 34.200 77.600 35.900 ;
        RECT 78.200 35.800 78.600 35.900 ;
        RECT 79.800 36.100 80.200 39.900 ;
        RECT 80.600 36.800 81.400 37.200 ;
        RECT 81.000 36.200 81.300 36.800 ;
        RECT 81.700 36.200 82.100 39.900 ;
        RECT 84.900 39.200 85.300 39.900 ;
        RECT 84.900 38.800 85.800 39.200 ;
        RECT 84.200 36.800 84.600 37.200 ;
        RECT 84.200 36.200 84.500 36.800 ;
        RECT 84.900 36.200 85.300 38.800 ;
        RECT 80.600 36.100 81.300 36.200 ;
        RECT 79.800 35.900 81.300 36.100 ;
        RECT 81.600 35.900 82.100 36.200 ;
        RECT 83.800 35.900 84.500 36.200 ;
        RECT 84.800 35.900 85.300 36.200 ;
        RECT 79.800 35.800 81.000 35.900 ;
        RECT 75.800 34.100 76.200 34.200 ;
        RECT 75.800 33.800 76.600 34.100 ;
        RECT 77.300 33.800 78.600 34.200 ;
        RECT 76.200 33.600 76.600 33.800 ;
        RECT 75.900 33.100 77.700 33.300 ;
        RECT 78.200 33.100 78.500 33.800 ;
        RECT 65.400 33.000 67.400 33.100 ;
        RECT 61.200 32.200 63.200 32.500 ;
        RECT 61.200 32.100 61.800 32.200 ;
        RECT 61.400 31.100 61.800 32.100 ;
        RECT 62.900 31.800 63.400 32.200 ;
        RECT 63.000 31.100 63.400 31.800 ;
        RECT 65.400 31.100 65.800 33.000 ;
        RECT 67.000 31.100 67.400 33.000 ;
        RECT 67.800 31.100 68.200 33.100 ;
        RECT 70.200 31.100 70.600 33.100 ;
        RECT 71.000 33.000 73.000 33.100 ;
        RECT 71.000 31.100 71.400 33.000 ;
        RECT 72.600 31.100 73.000 33.000 ;
        RECT 73.700 32.800 74.600 33.100 ;
        RECT 75.800 33.000 77.800 33.100 ;
        RECT 73.700 32.200 74.100 32.800 ;
        RECT 73.700 31.800 74.600 32.200 ;
        RECT 73.700 31.100 74.100 31.800 ;
        RECT 75.800 31.100 76.200 33.000 ;
        RECT 77.400 31.100 77.800 33.000 ;
        RECT 78.200 31.100 78.600 33.100 ;
        RECT 79.000 32.400 79.400 33.200 ;
        RECT 79.800 31.100 80.200 35.800 ;
        RECT 81.600 35.200 81.900 35.900 ;
        RECT 83.800 35.800 84.200 35.900 ;
        RECT 81.400 34.800 81.900 35.200 ;
        RECT 81.600 34.200 81.900 34.800 ;
        RECT 82.200 34.400 82.600 35.200 ;
        RECT 84.800 34.200 85.100 35.900 ;
        RECT 85.400 35.100 85.800 35.200 ;
        RECT 86.200 35.100 86.600 35.200 ;
        RECT 85.400 34.800 86.600 35.100 ;
        RECT 85.400 34.400 85.800 34.800 ;
        RECT 80.600 33.800 81.900 34.200 ;
        RECT 83.000 34.100 83.400 34.200 ;
        RECT 82.600 33.800 83.400 34.100 ;
        RECT 83.800 33.800 85.100 34.200 ;
        RECT 86.200 34.100 86.600 34.200 ;
        RECT 85.800 33.800 86.600 34.100 ;
        RECT 80.700 33.100 81.000 33.800 ;
        RECT 82.600 33.600 83.000 33.800 ;
        RECT 81.500 33.100 83.300 33.300 ;
        RECT 83.900 33.100 84.200 33.800 ;
        RECT 85.800 33.600 86.200 33.800 ;
        RECT 84.700 33.100 86.500 33.300 ;
        RECT 80.600 31.100 81.000 33.100 ;
        RECT 81.400 33.000 83.400 33.100 ;
        RECT 81.400 31.100 81.800 33.000 ;
        RECT 83.000 31.100 83.400 33.000 ;
        RECT 83.800 31.100 84.200 33.100 ;
        RECT 84.600 33.000 86.600 33.100 ;
        RECT 84.600 31.100 85.000 33.000 ;
        RECT 86.200 31.100 86.600 33.000 ;
        RECT 87.000 31.100 87.400 39.900 ;
        RECT 89.900 36.200 90.300 39.900 ;
        RECT 90.600 36.800 91.000 37.200 ;
        RECT 90.700 36.200 91.000 36.800 ;
        RECT 89.900 35.900 90.400 36.200 ;
        RECT 90.700 35.900 91.400 36.200 ;
        RECT 90.100 35.200 90.400 35.900 ;
        RECT 91.000 35.800 91.400 35.900 ;
        RECT 92.600 36.100 93.000 39.900 ;
        RECT 93.400 36.100 93.800 36.600 ;
        RECT 92.600 35.800 93.800 36.100 ;
        RECT 94.200 36.100 94.600 39.900 ;
        RECT 95.000 36.100 95.400 36.200 ;
        RECT 94.200 35.800 95.400 36.100 ;
        RECT 89.400 34.400 89.800 35.200 ;
        RECT 90.100 34.800 90.600 35.200 ;
        RECT 90.100 34.200 90.400 34.800 ;
        RECT 87.800 33.400 88.200 34.200 ;
        RECT 88.600 34.100 89.000 34.200 ;
        RECT 88.600 33.800 89.400 34.100 ;
        RECT 90.100 33.800 91.400 34.200 ;
        RECT 89.000 33.600 89.400 33.800 ;
        RECT 88.700 33.100 90.500 33.300 ;
        RECT 91.000 33.100 91.300 33.800 ;
        RECT 88.600 33.000 90.600 33.100 ;
        RECT 88.600 31.100 89.000 33.000 ;
        RECT 90.200 31.100 90.600 33.000 ;
        RECT 91.000 31.100 91.400 33.100 ;
        RECT 92.600 31.100 93.000 35.800 ;
        RECT 94.200 33.100 94.600 35.800 ;
        RECT 93.700 32.800 94.600 33.100 ;
        RECT 93.700 31.100 94.100 32.800 ;
        RECT 2.200 27.600 2.600 29.900 ;
        RECT 3.300 28.200 3.700 29.900 ;
        RECT 3.300 27.900 4.200 28.200 ;
        RECT 1.500 27.300 2.600 27.600 ;
        RECT 1.500 25.800 1.800 27.300 ;
        RECT 2.200 26.100 2.600 26.600 ;
        RECT 3.800 26.100 4.200 27.900 ;
        RECT 4.600 26.800 5.000 27.600 ;
        RECT 6.000 27.100 6.400 29.900 ;
        RECT 8.600 27.900 9.000 29.900 ;
        RECT 9.400 28.000 9.800 29.900 ;
        RECT 11.000 28.000 11.400 29.900 ;
        RECT 14.200 28.900 14.600 29.900 ;
        RECT 15.800 29.200 16.200 29.900 ;
        RECT 9.400 27.900 11.400 28.000 ;
        RECT 14.000 28.800 14.600 28.900 ;
        RECT 15.700 28.800 16.200 29.200 ;
        RECT 14.000 28.500 16.000 28.800 ;
        RECT 8.700 27.200 9.000 27.900 ;
        RECT 9.500 27.700 11.300 27.900 ;
        RECT 10.600 27.200 11.000 27.400 ;
        RECT 5.500 26.900 6.400 27.100 ;
        RECT 5.500 26.800 6.300 26.900 ;
        RECT 8.600 26.800 9.900 27.200 ;
        RECT 10.600 27.100 11.400 27.200 ;
        RECT 11.800 27.100 12.200 27.200 ;
        RECT 10.600 26.900 12.200 27.100 ;
        RECT 11.000 26.800 12.200 26.900 ;
        RECT 2.200 25.800 4.200 26.100 ;
        RECT 1.200 25.400 1.800 25.800 ;
        RECT 1.500 25.100 1.800 25.400 ;
        RECT 1.500 24.800 2.600 25.100 ;
        RECT 2.200 21.100 2.600 24.800 ;
        RECT 3.000 24.400 3.400 25.200 ;
        RECT 3.800 21.100 4.200 25.800 ;
        RECT 5.500 25.200 5.800 26.800 ;
        RECT 6.200 25.800 7.400 26.200 ;
        RECT 9.600 26.100 9.900 26.800 ;
        RECT 7.800 25.800 9.900 26.100 ;
        RECT 10.200 25.800 10.600 26.600 ;
        RECT 5.400 24.800 5.800 25.200 ;
        RECT 7.800 24.800 8.200 25.800 ;
        RECT 8.600 25.100 9.000 25.200 ;
        RECT 9.600 25.100 9.900 25.800 ;
        RECT 14.000 25.200 14.300 28.500 ;
        RECT 15.800 27.800 17.000 28.200 ;
        RECT 18.200 27.900 18.600 29.900 ;
        RECT 19.000 28.000 19.400 29.900 ;
        RECT 20.600 28.000 21.000 29.900 ;
        RECT 19.000 27.900 21.000 28.000 ;
        RECT 21.400 27.900 21.800 29.900 ;
        RECT 22.200 28.000 22.600 29.900 ;
        RECT 23.800 28.000 24.200 29.900 ;
        RECT 25.400 28.900 25.800 29.900 ;
        RECT 22.200 27.900 24.200 28.000 ;
        RECT 18.300 27.200 18.600 27.900 ;
        RECT 19.100 27.700 20.900 27.900 ;
        RECT 20.200 27.200 20.600 27.400 ;
        RECT 21.500 27.200 21.800 27.900 ;
        RECT 22.300 27.700 24.100 27.900 ;
        RECT 24.600 27.800 25.000 28.600 ;
        RECT 25.500 27.800 25.800 28.900 ;
        RECT 27.000 27.900 27.400 29.900 ;
        RECT 25.500 27.500 26.700 27.800 ;
        RECT 23.400 27.200 23.800 27.400 ;
        RECT 15.400 27.100 16.200 27.200 ;
        RECT 16.600 27.100 17.000 27.200 ;
        RECT 15.400 26.800 17.000 27.100 ;
        RECT 18.200 26.800 19.500 27.200 ;
        RECT 20.200 26.900 21.000 27.200 ;
        RECT 20.600 26.800 21.000 26.900 ;
        RECT 21.400 26.800 22.700 27.200 ;
        RECT 23.400 26.900 24.200 27.200 ;
        RECT 23.800 26.800 24.200 26.900 ;
        RECT 14.600 25.800 15.400 26.200 ;
        RECT 8.600 24.800 9.300 25.100 ;
        RECT 9.600 24.800 10.100 25.100 ;
        RECT 12.600 24.900 14.300 25.200 ;
        RECT 18.200 25.100 18.600 25.200 ;
        RECT 19.200 25.100 19.500 26.800 ;
        RECT 19.800 25.800 20.200 26.600 ;
        RECT 21.400 25.100 21.800 25.200 ;
        RECT 22.400 25.100 22.700 26.800 ;
        RECT 23.000 25.800 23.400 26.600 ;
        RECT 26.400 26.000 26.700 27.500 ;
        RECT 27.100 26.200 27.400 27.900 ;
        RECT 30.200 28.900 30.600 29.900 ;
        RECT 33.600 29.200 34.000 29.900 ;
        RECT 30.200 27.200 30.500 28.900 ;
        RECT 33.400 28.800 34.000 29.200 ;
        RECT 31.000 27.800 31.400 28.600 ;
        RECT 30.200 26.800 30.600 27.200 ;
        RECT 33.600 27.100 34.000 28.800 ;
        RECT 35.000 28.000 35.400 29.900 ;
        RECT 36.600 28.000 37.000 29.900 ;
        RECT 35.000 27.900 37.000 28.000 ;
        RECT 37.400 27.900 37.800 29.900 ;
        RECT 35.100 27.700 36.900 27.900 ;
        RECT 35.400 27.200 35.800 27.400 ;
        RECT 37.400 27.200 37.700 27.900 ;
        RECT 33.600 26.900 34.500 27.100 ;
        RECT 33.700 26.800 34.500 26.900 ;
        RECT 35.000 26.900 35.800 27.200 ;
        RECT 35.000 26.800 35.400 26.900 ;
        RECT 36.500 26.800 37.800 27.200 ;
        RECT 26.300 25.700 26.700 26.000 ;
        RECT 27.000 25.800 27.400 26.200 ;
        RECT 24.600 25.600 26.700 25.700 ;
        RECT 24.600 25.400 26.600 25.600 ;
        RECT 12.600 24.800 13.000 24.900 ;
        RECT 18.200 24.800 18.900 25.100 ;
        RECT 19.200 24.800 19.700 25.100 ;
        RECT 21.400 24.800 22.100 25.100 ;
        RECT 22.400 24.800 22.900 25.100 ;
        RECT 5.500 23.500 5.800 24.800 ;
        RECT 6.200 23.800 6.600 24.600 ;
        RECT 9.000 24.200 9.300 24.800 ;
        RECT 9.000 23.800 9.400 24.200 ;
        RECT 5.500 23.200 7.300 23.500 ;
        RECT 5.500 23.100 5.800 23.200 ;
        RECT 5.400 21.100 5.800 23.100 ;
        RECT 7.000 23.100 7.300 23.200 ;
        RECT 7.000 21.100 7.400 23.100 ;
        RECT 9.700 21.100 10.100 24.800 ;
        RECT 12.700 24.500 13.000 24.800 ;
        RECT 13.500 24.500 15.300 24.600 ;
        RECT 11.800 21.500 12.200 24.500 ;
        RECT 12.600 21.700 13.000 24.500 ;
        RECT 13.400 24.300 15.300 24.500 ;
        RECT 11.900 21.400 12.200 21.500 ;
        RECT 13.400 21.500 13.800 24.300 ;
        RECT 15.000 24.100 15.300 24.300 ;
        RECT 15.900 24.400 17.700 24.700 ;
        RECT 15.900 24.100 16.200 24.400 ;
        RECT 13.400 21.400 13.700 21.500 ;
        RECT 11.900 21.100 13.700 21.400 ;
        RECT 14.200 21.400 14.600 24.000 ;
        RECT 15.000 21.700 15.400 24.100 ;
        RECT 15.800 21.400 16.200 24.100 ;
        RECT 14.200 21.100 16.200 21.400 ;
        RECT 17.400 24.100 17.700 24.400 ;
        RECT 18.600 24.200 18.900 24.800 ;
        RECT 17.400 21.100 17.800 24.100 ;
        RECT 18.600 23.800 19.000 24.200 ;
        RECT 19.300 21.100 19.700 24.800 ;
        RECT 21.800 24.200 22.100 24.800 ;
        RECT 21.800 23.800 22.200 24.200 ;
        RECT 22.500 23.200 22.900 24.800 ;
        RECT 22.500 22.800 23.400 23.200 ;
        RECT 22.500 21.100 22.900 22.800 ;
        RECT 24.600 21.100 25.000 25.400 ;
        RECT 27.100 25.200 27.400 25.800 ;
        RECT 29.400 25.400 29.800 26.200 ;
        RECT 27.000 25.100 27.400 25.200 ;
        RECT 30.200 25.100 30.500 26.800 ;
        RECT 32.600 25.800 33.800 26.200 ;
        RECT 31.800 25.100 32.200 25.600 ;
        RECT 34.200 25.200 34.500 26.800 ;
        RECT 35.800 25.800 36.200 26.600 ;
        RECT 26.700 24.800 27.400 25.100 ;
        RECT 26.700 21.100 27.100 24.800 ;
        RECT 29.700 24.700 30.600 25.100 ;
        RECT 31.800 24.800 32.900 25.100 ;
        RECT 28.600 24.100 29.000 24.200 ;
        RECT 29.700 24.100 30.100 24.700 ;
        RECT 28.600 23.800 30.100 24.100 ;
        RECT 32.600 24.200 32.900 24.800 ;
        RECT 34.200 24.800 34.600 25.200 ;
        RECT 36.500 25.100 36.800 26.800 ;
        RECT 37.400 25.100 37.800 25.200 ;
        RECT 38.200 25.100 38.600 29.900 ;
        RECT 40.600 28.900 41.000 29.900 ;
        RECT 39.000 27.800 39.400 28.600 ;
        RECT 39.000 27.100 39.300 27.800 ;
        RECT 40.700 27.200 41.000 28.900 ;
        RECT 42.200 28.000 42.600 29.900 ;
        RECT 43.800 28.000 44.200 29.900 ;
        RECT 42.200 27.900 44.200 28.000 ;
        RECT 44.600 27.900 45.000 29.900 ;
        RECT 42.300 27.700 44.100 27.900 ;
        RECT 42.600 27.200 43.000 27.400 ;
        RECT 44.600 27.200 44.900 27.900 ;
        RECT 40.600 27.100 41.000 27.200 ;
        RECT 39.000 26.800 41.000 27.100 ;
        RECT 42.200 26.900 43.000 27.200 ;
        RECT 42.200 26.800 42.600 26.900 ;
        RECT 43.700 26.800 45.000 27.200 ;
        RECT 40.700 25.100 41.000 26.800 ;
        RECT 41.400 25.400 41.800 26.200 ;
        RECT 43.000 25.800 43.400 26.600 ;
        RECT 43.700 26.200 44.000 26.800 ;
        RECT 43.700 25.800 44.200 26.200 ;
        RECT 44.600 26.100 45.000 26.200 ;
        RECT 45.400 26.100 45.800 29.900 ;
        RECT 48.500 27.900 49.300 29.900 ;
        RECT 47.800 26.400 48.200 27.200 ;
        RECT 48.700 26.200 49.000 27.900 ;
        RECT 51.000 27.800 51.400 28.600 ;
        RECT 49.400 26.800 49.800 27.200 ;
        RECT 49.400 26.600 49.700 26.800 ;
        RECT 49.300 26.200 49.700 26.600 ;
        RECT 47.000 26.100 47.400 26.200 ;
        RECT 44.600 25.800 47.800 26.100 ;
        RECT 48.600 25.800 49.000 26.200 ;
        RECT 43.700 25.100 44.000 25.800 ;
        RECT 44.600 25.100 45.000 25.200 ;
        RECT 36.300 24.800 36.800 25.100 ;
        RECT 37.100 24.800 38.600 25.100 ;
        RECT 32.600 23.800 33.000 24.200 ;
        RECT 33.400 23.800 33.800 24.600 ;
        RECT 29.700 21.100 30.100 23.800 ;
        RECT 34.200 23.500 34.500 24.800 ;
        RECT 32.700 23.200 34.500 23.500 ;
        RECT 32.700 23.100 33.000 23.200 ;
        RECT 32.600 21.100 33.000 23.100 ;
        RECT 34.200 23.100 34.500 23.200 ;
        RECT 34.200 21.100 34.600 23.100 ;
        RECT 36.300 21.100 36.700 24.800 ;
        RECT 37.100 24.200 37.400 24.800 ;
        RECT 37.000 23.800 37.400 24.200 ;
        RECT 38.200 21.100 38.600 24.800 ;
        RECT 40.600 24.700 41.500 25.100 ;
        RECT 41.100 21.100 41.500 24.700 ;
        RECT 43.500 24.800 44.000 25.100 ;
        RECT 44.300 24.800 45.000 25.100 ;
        RECT 43.500 21.100 43.900 24.800 ;
        RECT 44.300 24.200 44.600 24.800 ;
        RECT 44.200 23.800 44.600 24.200 ;
        RECT 45.400 21.100 45.800 25.800 ;
        RECT 47.400 25.600 47.800 25.800 ;
        RECT 48.700 25.700 49.000 25.800 ;
        RECT 48.700 25.400 49.700 25.700 ;
        RECT 50.200 25.400 50.600 26.200 ;
        RECT 51.000 26.100 51.400 26.200 ;
        RECT 51.800 26.100 52.200 29.900 ;
        RECT 53.900 27.900 54.700 29.900 ;
        RECT 58.200 27.900 58.600 29.900 ;
        RECT 58.900 28.200 59.300 28.600 ;
        RECT 53.400 26.800 53.800 27.200 ;
        RECT 53.500 26.600 53.800 26.800 ;
        RECT 53.500 26.200 53.900 26.600 ;
        RECT 54.200 26.200 54.500 27.900 ;
        RECT 55.000 26.400 55.400 27.200 ;
        RECT 57.400 26.400 57.800 27.200 ;
        RECT 51.000 25.800 52.200 26.100 ;
        RECT 49.400 25.100 49.700 25.400 ;
        RECT 47.000 24.800 49.000 25.100 ;
        RECT 47.000 21.100 47.400 24.800 ;
        RECT 48.600 21.400 49.000 24.800 ;
        RECT 49.400 21.700 49.800 25.100 ;
        RECT 50.200 21.400 50.600 25.100 ;
        RECT 48.600 21.100 50.600 21.400 ;
        RECT 51.800 21.100 52.200 25.800 ;
        RECT 54.200 25.800 54.600 26.200 ;
        RECT 55.800 26.100 56.200 26.200 ;
        RECT 55.400 25.800 56.200 26.100 ;
        RECT 56.600 26.100 57.000 26.200 ;
        RECT 58.200 26.100 58.500 27.900 ;
        RECT 59.000 27.800 59.400 28.200 ;
        RECT 61.400 27.900 61.800 29.900 ;
        RECT 62.100 28.200 62.500 28.600 ;
        RECT 60.600 26.400 61.000 27.200 ;
        RECT 59.000 26.100 59.400 26.200 ;
        RECT 56.600 25.800 57.400 26.100 ;
        RECT 58.200 25.800 59.400 26.100 ;
        RECT 59.800 26.100 60.200 26.200 ;
        RECT 61.400 26.100 61.700 27.900 ;
        RECT 62.200 27.800 62.600 28.200 ;
        RECT 63.000 28.000 63.400 29.900 ;
        RECT 64.600 28.000 65.000 29.900 ;
        RECT 63.000 27.900 65.000 28.000 ;
        RECT 65.400 27.900 65.800 29.900 ;
        RECT 67.000 28.900 67.400 29.900 ;
        RECT 63.100 27.700 64.900 27.900 ;
        RECT 63.400 27.200 63.800 27.400 ;
        RECT 65.400 27.200 65.700 27.900 ;
        RECT 67.000 27.200 67.300 28.900 ;
        RECT 67.800 28.100 68.200 28.600 ;
        RECT 70.200 28.100 70.600 29.900 ;
        RECT 67.800 27.800 70.600 28.100 ;
        RECT 71.000 28.000 71.400 29.900 ;
        RECT 72.600 28.000 73.000 29.900 ;
        RECT 73.700 29.200 74.100 29.900 ;
        RECT 73.400 28.800 74.100 29.200 ;
        RECT 71.000 27.900 73.000 28.000 ;
        RECT 73.700 28.200 74.100 28.800 ;
        RECT 73.700 27.900 74.600 28.200 ;
        RECT 75.800 27.900 76.200 29.900 ;
        RECT 76.600 28.000 77.000 29.900 ;
        RECT 78.200 28.000 78.600 29.900 ;
        RECT 76.600 27.900 78.600 28.000 ;
        RECT 79.800 28.800 80.200 29.900 ;
        RECT 70.300 27.200 70.600 27.800 ;
        RECT 71.100 27.700 72.900 27.900 ;
        RECT 72.200 27.200 72.600 27.400 ;
        RECT 62.200 27.100 62.600 27.200 ;
        RECT 63.000 27.100 63.800 27.200 ;
        RECT 62.200 26.900 63.800 27.100 ;
        RECT 62.200 26.800 63.400 26.900 ;
        RECT 64.500 26.800 65.800 27.200 ;
        RECT 67.000 26.800 67.400 27.200 ;
        RECT 70.200 26.800 71.500 27.200 ;
        RECT 72.200 26.900 73.000 27.200 ;
        RECT 72.600 26.800 73.000 26.900 ;
        RECT 62.200 26.100 62.600 26.200 ;
        RECT 59.800 25.800 60.600 26.100 ;
        RECT 61.400 25.800 62.600 26.100 ;
        RECT 63.800 25.800 64.200 26.600 ;
        RECT 64.500 26.100 64.800 26.800 ;
        RECT 66.200 26.100 66.600 26.200 ;
        RECT 64.500 25.800 66.600 26.100 ;
        RECT 54.200 25.700 54.500 25.800 ;
        RECT 53.500 25.400 54.500 25.700 ;
        RECT 55.400 25.600 55.800 25.800 ;
        RECT 57.000 25.600 57.400 25.800 ;
        RECT 53.500 25.100 53.800 25.400 ;
        RECT 59.000 25.100 59.300 25.800 ;
        RECT 60.200 25.600 60.600 25.800 ;
        RECT 62.200 25.100 62.500 25.800 ;
        RECT 64.500 25.100 64.800 25.800 ;
        RECT 66.200 25.400 66.600 25.800 ;
        RECT 65.400 25.100 65.800 25.200 ;
        RECT 67.000 25.100 67.300 26.800 ;
        RECT 70.200 25.100 70.600 25.200 ;
        RECT 71.200 25.100 71.500 26.800 ;
        RECT 71.800 25.800 72.200 26.600 ;
        RECT 52.600 21.400 53.000 25.100 ;
        RECT 53.400 21.700 53.800 25.100 ;
        RECT 54.200 24.800 56.200 25.100 ;
        RECT 54.200 21.400 54.600 24.800 ;
        RECT 52.600 21.100 54.600 21.400 ;
        RECT 55.800 21.100 56.200 24.800 ;
        RECT 56.600 24.800 58.600 25.100 ;
        RECT 56.600 21.100 57.000 24.800 ;
        RECT 58.200 21.100 58.600 24.800 ;
        RECT 59.000 21.100 59.400 25.100 ;
        RECT 59.800 24.800 61.800 25.100 ;
        RECT 59.800 21.100 60.200 24.800 ;
        RECT 61.400 21.100 61.800 24.800 ;
        RECT 62.200 21.100 62.600 25.100 ;
        RECT 64.300 24.800 64.800 25.100 ;
        RECT 65.100 24.800 65.800 25.100 ;
        RECT 64.300 21.100 64.700 24.800 ;
        RECT 65.100 24.200 65.400 24.800 ;
        RECT 65.000 23.800 65.400 24.200 ;
        RECT 66.500 24.700 67.400 25.100 ;
        RECT 70.200 24.800 70.900 25.100 ;
        RECT 71.200 24.800 71.700 25.100 ;
        RECT 66.500 22.200 66.900 24.700 ;
        RECT 70.600 24.200 70.900 24.800 ;
        RECT 70.600 23.800 71.000 24.200 ;
        RECT 66.200 21.800 66.900 22.200 ;
        RECT 66.500 21.100 66.900 21.800 ;
        RECT 71.300 21.100 71.700 24.800 ;
        RECT 73.400 24.400 73.800 25.200 ;
        RECT 74.200 21.100 74.600 27.900 ;
        RECT 75.000 26.800 75.400 27.600 ;
        RECT 75.900 27.200 76.200 27.900 ;
        RECT 76.700 27.700 78.500 27.900 ;
        RECT 77.800 27.200 78.200 27.400 ;
        RECT 79.800 27.200 80.100 28.800 ;
        RECT 80.600 27.800 81.000 28.600 ;
        RECT 83.000 27.900 83.400 29.900 ;
        RECT 83.700 28.200 84.100 28.600 ;
        RECT 75.800 26.800 77.100 27.200 ;
        RECT 77.800 27.100 78.600 27.200 ;
        RECT 79.000 27.100 79.400 27.200 ;
        RECT 77.800 26.900 79.400 27.100 ;
        RECT 78.200 26.800 79.400 26.900 ;
        RECT 79.800 26.800 80.200 27.200 ;
        RECT 80.600 27.100 80.900 27.800 ;
        RECT 82.200 27.100 82.600 27.200 ;
        RECT 80.600 26.800 82.600 27.100 ;
        RECT 75.800 25.100 76.200 25.200 ;
        RECT 76.800 25.100 77.100 26.800 ;
        RECT 77.400 25.800 77.800 26.600 ;
        RECT 78.200 26.100 78.600 26.200 ;
        RECT 79.000 26.100 79.400 26.200 ;
        RECT 78.200 25.800 79.400 26.100 ;
        RECT 79.000 25.400 79.400 25.800 ;
        RECT 79.800 25.100 80.100 26.800 ;
        RECT 82.200 26.400 82.600 26.800 ;
        RECT 80.600 26.100 81.000 26.200 ;
        RECT 81.400 26.100 81.800 26.200 ;
        RECT 83.000 26.100 83.300 27.900 ;
        RECT 83.800 27.800 84.200 28.200 ;
        RECT 84.600 27.900 85.000 29.900 ;
        RECT 85.400 28.000 85.800 29.900 ;
        RECT 87.000 28.000 87.400 29.900 ;
        RECT 85.400 27.900 87.400 28.000 ;
        RECT 84.700 27.200 85.000 27.900 ;
        RECT 85.500 27.700 87.300 27.900 ;
        RECT 86.600 27.200 87.000 27.400 ;
        RECT 83.800 27.100 84.200 27.200 ;
        RECT 84.600 27.100 85.900 27.200 ;
        RECT 83.800 26.800 85.900 27.100 ;
        RECT 86.600 26.900 87.400 27.200 ;
        RECT 87.000 26.800 87.400 26.900 ;
        RECT 83.800 26.100 84.200 26.200 ;
        RECT 80.600 25.800 82.200 26.100 ;
        RECT 83.000 25.800 84.200 26.100 ;
        RECT 81.800 25.600 82.200 25.800 ;
        RECT 83.800 25.100 84.100 25.800 ;
        RECT 84.600 25.100 85.000 25.200 ;
        RECT 85.600 25.100 85.900 26.800 ;
        RECT 86.200 25.800 86.600 26.600 ;
        RECT 75.800 24.800 76.500 25.100 ;
        RECT 76.800 24.800 77.300 25.100 ;
        RECT 76.200 24.200 76.500 24.800 ;
        RECT 76.200 23.800 76.600 24.200 ;
        RECT 76.900 21.100 77.300 24.800 ;
        RECT 79.300 24.700 80.200 25.100 ;
        RECT 81.400 24.800 83.400 25.100 ;
        RECT 79.300 21.100 79.700 24.700 ;
        RECT 81.400 21.100 81.800 24.800 ;
        RECT 83.000 21.100 83.400 24.800 ;
        RECT 83.800 24.800 85.300 25.100 ;
        RECT 85.600 24.800 86.100 25.100 ;
        RECT 83.800 21.100 84.200 24.800 ;
        RECT 85.000 24.200 85.300 24.800 ;
        RECT 85.000 23.800 85.400 24.200 ;
        RECT 85.700 21.100 86.100 24.800 ;
        RECT 87.800 21.100 88.200 29.900 ;
        RECT 89.700 28.200 90.100 29.900 ;
        RECT 92.600 28.900 93.000 29.900 ;
        RECT 89.400 27.800 90.600 28.200 ;
        RECT 88.600 26.800 89.000 27.600 ;
        RECT 89.400 27.200 89.700 27.800 ;
        RECT 89.400 26.800 89.800 27.200 ;
        RECT 89.400 24.400 89.800 25.200 ;
        RECT 90.200 21.100 90.600 27.800 ;
        RECT 91.000 26.800 91.400 27.600 ;
        RECT 92.600 27.200 92.900 28.900 ;
        RECT 93.400 28.100 93.800 28.600 ;
        RECT 94.200 28.100 94.600 29.900 ;
        RECT 93.400 27.800 94.600 28.100 ;
        RECT 95.000 28.000 95.400 29.900 ;
        RECT 96.600 28.000 97.000 29.900 ;
        RECT 95.000 27.900 97.000 28.000 ;
        RECT 94.300 27.200 94.600 27.800 ;
        RECT 95.100 27.700 96.900 27.900 ;
        RECT 96.200 27.200 96.600 27.400 ;
        RECT 92.600 26.800 93.000 27.200 ;
        RECT 94.200 26.800 95.500 27.200 ;
        RECT 96.200 26.900 97.000 27.200 ;
        RECT 96.600 26.800 97.000 26.900 ;
        RECT 91.800 25.400 92.200 26.200 ;
        RECT 92.600 25.100 92.900 26.800 ;
        RECT 94.200 25.100 94.600 25.200 ;
        RECT 95.200 25.100 95.500 26.800 ;
        RECT 95.800 25.800 96.200 26.600 ;
        RECT 92.100 24.700 93.000 25.100 ;
        RECT 94.200 24.800 94.900 25.100 ;
        RECT 95.200 24.800 95.700 25.100 ;
        RECT 92.100 22.200 92.500 24.700 ;
        RECT 94.600 24.200 94.900 24.800 ;
        RECT 94.600 23.800 95.000 24.200 ;
        RECT 92.100 21.800 93.000 22.200 ;
        RECT 92.100 21.100 92.500 21.800 ;
        RECT 95.300 21.100 95.700 24.800 ;
        RECT 0.700 19.600 2.500 19.900 ;
        RECT 0.700 19.500 1.000 19.600 ;
        RECT 0.600 16.500 1.000 19.500 ;
        RECT 2.200 19.500 2.500 19.600 ;
        RECT 3.000 19.600 5.000 19.900 ;
        RECT 1.400 16.500 1.800 19.300 ;
        RECT 2.200 16.700 2.600 19.500 ;
        RECT 3.000 17.000 3.400 19.600 ;
        RECT 3.800 16.900 4.200 19.300 ;
        RECT 4.600 16.900 5.000 19.600 ;
        RECT 3.800 16.700 4.100 16.900 ;
        RECT 2.200 16.500 4.100 16.700 ;
        RECT 1.500 16.200 1.800 16.500 ;
        RECT 2.300 16.400 4.100 16.500 ;
        RECT 4.700 16.600 5.000 16.900 ;
        RECT 6.200 16.900 6.600 19.900 ;
        RECT 8.300 17.200 8.700 19.900 ;
        RECT 10.200 17.900 10.600 19.900 ;
        RECT 10.300 17.800 10.600 17.900 ;
        RECT 11.800 17.900 12.200 19.900 ;
        RECT 11.800 17.800 12.100 17.900 ;
        RECT 10.300 17.500 12.100 17.800 ;
        RECT 6.200 16.600 6.500 16.900 ;
        RECT 7.800 16.800 8.700 17.200 ;
        RECT 9.000 16.800 9.800 17.200 ;
        RECT 4.700 16.300 6.500 16.600 ;
        RECT 1.400 16.100 1.800 16.200 ;
        RECT 8.300 16.200 8.700 16.800 ;
        RECT 9.100 16.200 9.400 16.800 ;
        RECT 10.300 16.200 10.600 17.500 ;
        RECT 11.000 16.400 11.400 17.200 ;
        RECT 1.400 15.800 3.100 16.100 ;
        RECT 8.300 15.900 8.800 16.200 ;
        RECT 9.100 15.900 9.800 16.200 ;
        RECT 2.800 14.200 3.100 15.800 ;
        RECT 3.400 14.800 4.200 15.200 ;
        RECT 8.500 14.200 8.800 15.900 ;
        RECT 9.400 15.800 9.800 15.900 ;
        RECT 10.200 15.800 10.600 16.200 ;
        RECT 9.400 15.100 9.800 15.200 ;
        RECT 10.300 15.100 10.600 15.800 ;
        RECT 12.600 15.400 13.000 16.200 ;
        RECT 13.400 15.800 13.800 16.200 ;
        RECT 9.400 14.800 10.600 15.100 ;
        RECT 11.400 14.800 12.200 15.200 ;
        RECT 13.400 15.100 13.700 15.800 ;
        RECT 14.200 15.100 14.600 19.900 ;
        RECT 15.000 15.800 15.400 17.200 ;
        RECT 15.800 15.800 16.200 16.600 ;
        RECT 13.400 14.800 14.600 15.100 ;
        RECT 15.000 15.100 15.400 15.200 ;
        RECT 16.600 15.100 17.000 19.900 ;
        RECT 18.200 16.200 18.600 19.900 ;
        RECT 19.800 16.200 20.200 19.900 ;
        RECT 18.200 15.900 20.200 16.200 ;
        RECT 20.600 15.900 21.000 19.900 ;
        RECT 21.800 16.800 22.200 17.200 ;
        RECT 21.800 16.200 22.100 16.800 ;
        RECT 22.500 16.200 22.900 19.900 ;
        RECT 21.400 15.900 22.100 16.200 ;
        RECT 22.400 15.900 22.900 16.200 ;
        RECT 18.600 15.200 19.000 15.400 ;
        RECT 20.600 15.200 20.900 15.900 ;
        RECT 21.400 15.800 21.800 15.900 ;
        RECT 21.400 15.200 21.700 15.800 ;
        RECT 15.000 14.800 17.000 15.100 ;
        RECT 18.200 14.900 19.000 15.200 ;
        RECT 19.800 14.900 21.000 15.200 ;
        RECT 18.200 14.800 18.600 14.900 ;
        RECT 10.300 14.200 10.600 14.800 ;
        RECT 2.800 13.800 3.400 14.200 ;
        RECT 4.200 13.800 5.000 14.200 ;
        RECT 8.500 13.800 9.800 14.200 ;
        RECT 10.300 14.100 11.100 14.200 ;
        RECT 10.300 13.900 11.200 14.100 ;
        RECT 2.800 12.500 3.100 13.800 ;
        RECT 4.900 12.800 5.800 13.200 ;
        RECT 7.100 13.100 8.900 13.300 ;
        RECT 9.400 13.100 9.700 13.800 ;
        RECT 7.000 13.000 9.000 13.100 ;
        RECT 2.800 12.200 4.800 12.500 ;
        RECT 2.800 12.100 3.400 12.200 ;
        RECT 3.000 11.100 3.400 12.100 ;
        RECT 4.500 12.100 4.800 12.200 ;
        RECT 4.500 11.800 5.000 12.100 ;
        RECT 4.600 11.100 5.000 11.800 ;
        RECT 7.000 11.100 7.400 13.000 ;
        RECT 8.600 11.100 9.000 13.000 ;
        RECT 9.400 11.100 9.800 13.100 ;
        RECT 10.800 11.100 11.200 13.900 ;
        RECT 13.400 13.400 13.800 14.200 ;
        RECT 14.200 13.100 14.600 14.800 ;
        RECT 16.600 13.100 17.000 14.800 ;
        RECT 19.000 13.800 19.400 14.600 ;
        RECT 14.200 12.800 15.100 13.100 ;
        RECT 14.700 11.100 15.100 12.800 ;
        RECT 16.100 12.800 17.000 13.100 ;
        RECT 19.800 13.200 20.100 14.900 ;
        RECT 20.600 14.800 21.000 14.900 ;
        RECT 21.400 14.800 21.800 15.200 ;
        RECT 22.400 14.200 22.700 15.900 ;
        RECT 23.000 14.400 23.400 15.200 ;
        RECT 21.400 13.800 22.700 14.200 ;
        RECT 23.800 14.100 24.200 14.200 ;
        RECT 23.400 13.800 24.200 14.100 ;
        RECT 16.100 11.100 16.500 12.800 ;
        RECT 19.800 11.100 20.200 13.200 ;
        RECT 20.600 13.100 21.000 13.200 ;
        RECT 21.500 13.100 21.800 13.800 ;
        RECT 23.400 13.600 23.800 13.800 ;
        RECT 22.300 13.100 24.100 13.300 ;
        RECT 25.400 13.100 25.800 19.900 ;
        RECT 28.600 13.400 29.000 14.200 ;
        RECT 29.400 14.100 29.800 19.900 ;
        RECT 31.800 17.900 32.200 19.900 ;
        RECT 31.900 17.800 32.200 17.900 ;
        RECT 33.400 17.900 33.800 19.900 ;
        RECT 33.400 17.800 33.700 17.900 ;
        RECT 31.900 17.500 33.700 17.800 ;
        RECT 32.600 17.100 33.000 17.200 ;
        RECT 30.200 16.800 33.000 17.100 ;
        RECT 30.200 15.800 30.600 16.800 ;
        RECT 32.600 16.400 33.000 16.800 ;
        RECT 33.400 16.200 33.700 17.500 ;
        RECT 35.500 16.200 35.900 19.900 ;
        RECT 36.200 16.800 36.600 17.200 ;
        RECT 36.300 16.200 36.600 16.800 ;
        RECT 38.700 16.300 39.100 19.900 ;
        RECT 31.000 15.400 31.400 16.200 ;
        RECT 33.400 15.800 33.800 16.200 ;
        RECT 35.500 15.900 36.000 16.200 ;
        RECT 36.300 15.900 37.000 16.200 ;
        RECT 38.200 15.900 39.100 16.300 ;
        RECT 39.800 15.900 40.200 19.900 ;
        RECT 40.600 16.200 41.000 19.900 ;
        RECT 42.200 16.200 42.600 19.900 ;
        RECT 40.600 15.900 42.600 16.200 ;
        RECT 43.000 16.200 43.400 19.900 ;
        RECT 44.600 16.200 45.000 19.900 ;
        RECT 43.000 15.900 45.000 16.200 ;
        RECT 45.400 15.900 45.800 19.900 ;
        RECT 46.200 17.900 46.600 19.900 ;
        RECT 46.300 17.800 46.600 17.900 ;
        RECT 47.800 17.900 48.200 19.900 ;
        RECT 49.400 19.600 51.400 19.900 ;
        RECT 47.800 17.800 48.100 17.900 ;
        RECT 46.300 17.500 48.100 17.800 ;
        RECT 46.300 16.200 46.600 17.500 ;
        RECT 47.000 16.400 47.400 17.200 ;
        RECT 30.200 14.800 30.600 15.200 ;
        RECT 31.800 14.800 32.600 15.200 ;
        RECT 30.200 14.100 30.500 14.800 ;
        RECT 33.400 14.200 33.700 15.800 ;
        RECT 34.200 15.100 34.600 15.200 ;
        RECT 35.000 15.100 35.400 15.200 ;
        RECT 34.200 14.800 35.400 15.100 ;
        RECT 35.000 14.400 35.400 14.800 ;
        RECT 35.700 14.200 36.000 15.900 ;
        RECT 36.600 15.800 37.000 15.900 ;
        RECT 38.300 14.200 38.600 15.900 ;
        RECT 39.000 14.800 39.400 15.600 ;
        RECT 39.900 15.200 40.200 15.900 ;
        RECT 41.800 15.200 42.200 15.400 ;
        RECT 43.400 15.200 43.800 15.400 ;
        RECT 45.400 15.200 45.700 15.900 ;
        RECT 46.200 15.800 46.600 16.200 ;
        RECT 39.800 14.900 41.000 15.200 ;
        RECT 41.800 14.900 42.600 15.200 ;
        RECT 39.800 14.800 40.200 14.900 ;
        RECT 32.900 14.100 33.700 14.200 ;
        RECT 29.400 13.800 30.500 14.100 ;
        RECT 32.800 13.900 33.700 14.100 ;
        RECT 34.200 14.100 34.600 14.200 ;
        RECT 29.400 13.100 29.800 13.800 ;
        RECT 20.600 12.800 21.800 13.100 ;
        RECT 20.500 12.400 20.900 12.800 ;
        RECT 21.400 11.100 21.800 12.800 ;
        RECT 22.200 13.000 24.200 13.100 ;
        RECT 22.200 11.100 22.600 13.000 ;
        RECT 23.800 11.100 24.200 13.000 ;
        RECT 25.400 12.800 26.300 13.100 ;
        RECT 29.400 12.800 30.300 13.100 ;
        RECT 25.900 12.200 26.300 12.800 ;
        RECT 25.900 11.800 26.600 12.200 ;
        RECT 25.900 11.100 26.300 11.800 ;
        RECT 29.900 11.100 30.300 12.800 ;
        RECT 32.800 11.100 33.200 13.900 ;
        RECT 34.200 13.800 35.000 14.100 ;
        RECT 35.700 13.800 37.000 14.200 ;
        RECT 38.200 13.800 38.600 14.200 ;
        RECT 34.600 13.600 35.000 13.800 ;
        RECT 34.300 13.100 36.100 13.300 ;
        RECT 36.600 13.100 36.900 13.800 ;
        RECT 34.200 13.000 36.200 13.100 ;
        RECT 34.200 11.100 34.600 13.000 ;
        RECT 35.800 11.100 36.200 13.000 ;
        RECT 36.600 11.100 37.000 13.100 ;
        RECT 37.400 12.400 37.800 13.200 ;
        RECT 38.300 13.100 38.600 13.800 ;
        RECT 39.000 13.800 39.400 14.200 ;
        RECT 39.000 13.100 39.300 13.800 ;
        RECT 38.200 12.800 39.300 13.100 ;
        RECT 39.800 12.800 40.200 13.200 ;
        RECT 40.700 13.100 41.000 14.900 ;
        RECT 42.200 14.800 42.600 14.900 ;
        RECT 43.000 14.900 43.800 15.200 ;
        RECT 44.600 14.900 45.800 15.200 ;
        RECT 43.000 14.800 43.400 14.900 ;
        RECT 44.600 14.800 45.000 14.900 ;
        RECT 45.400 14.800 45.800 14.900 ;
        RECT 41.400 13.800 41.800 14.600 ;
        RECT 43.800 13.800 44.200 14.600 ;
        RECT 38.300 12.100 38.600 12.800 ;
        RECT 39.900 12.400 40.300 12.800 ;
        RECT 38.200 11.100 38.600 12.100 ;
        RECT 40.600 11.100 41.000 13.100 ;
        RECT 44.600 13.100 44.900 14.800 ;
        RECT 46.300 14.200 46.600 15.800 ;
        RECT 48.600 15.400 49.000 16.200 ;
        RECT 49.400 15.900 49.800 19.600 ;
        RECT 50.200 15.800 50.600 19.300 ;
        RECT 51.000 16.200 51.400 19.600 ;
        RECT 52.600 16.200 53.000 19.900 ;
        RECT 51.000 15.900 53.000 16.200 ;
        RECT 54.700 16.200 55.100 19.900 ;
        RECT 55.400 16.800 55.800 17.200 ;
        RECT 56.600 16.900 57.000 19.900 ;
        RECT 55.500 16.200 55.800 16.800 ;
        RECT 56.700 16.600 57.000 16.900 ;
        RECT 58.200 19.600 60.200 19.900 ;
        RECT 58.200 16.900 58.600 19.600 ;
        RECT 59.000 16.900 59.400 19.300 ;
        RECT 59.800 17.000 60.200 19.600 ;
        RECT 60.700 19.600 62.500 19.900 ;
        RECT 60.700 19.500 61.000 19.600 ;
        RECT 58.200 16.600 58.500 16.900 ;
        RECT 56.700 16.300 58.500 16.600 ;
        RECT 59.100 16.700 59.400 16.900 ;
        RECT 60.600 16.700 61.000 19.500 ;
        RECT 62.200 19.500 62.500 19.600 ;
        RECT 59.100 16.500 61.000 16.700 ;
        RECT 61.400 16.500 61.800 19.300 ;
        RECT 62.200 16.500 62.600 19.500 ;
        RECT 59.100 16.400 60.900 16.500 ;
        RECT 61.400 16.200 61.700 16.500 ;
        RECT 64.300 16.200 64.700 19.900 ;
        RECT 65.000 16.800 65.400 17.200 ;
        RECT 65.100 16.200 65.400 16.800 ;
        RECT 66.600 16.800 67.000 17.200 ;
        RECT 66.600 16.200 66.900 16.800 ;
        RECT 67.300 16.200 67.700 19.900 ;
        RECT 54.700 15.900 55.200 16.200 ;
        RECT 55.500 15.900 56.200 16.200 ;
        RECT 61.400 16.100 61.800 16.200 ;
        RECT 50.300 15.600 50.600 15.800 ;
        RECT 50.300 15.300 51.300 15.600 ;
        RECT 51.000 15.200 51.300 15.300 ;
        RECT 52.200 15.200 52.600 15.400 ;
        RECT 47.400 14.800 48.200 15.200 ;
        RECT 51.000 14.800 51.400 15.200 ;
        RECT 52.200 14.900 53.000 15.200 ;
        RECT 52.600 14.800 53.000 14.900 ;
        RECT 50.300 14.400 50.700 14.800 ;
        RECT 50.300 14.200 50.600 14.400 ;
        RECT 46.300 14.100 47.100 14.200 ;
        RECT 46.300 13.900 47.200 14.100 ;
        RECT 45.400 13.100 45.800 13.200 ;
        RECT 46.800 13.100 47.200 13.900 ;
        RECT 50.200 13.800 50.600 14.200 ;
        RECT 51.000 13.100 51.300 14.800 ;
        RECT 54.200 14.400 54.600 15.200 ;
        RECT 54.900 14.200 55.200 15.900 ;
        RECT 55.800 15.800 56.200 15.900 ;
        RECT 60.100 15.800 61.800 16.100 ;
        RECT 64.300 15.900 64.800 16.200 ;
        RECT 65.100 15.900 65.800 16.200 ;
        RECT 59.000 14.800 59.800 15.200 ;
        RECT 53.400 14.100 53.800 14.200 ;
        RECT 54.900 14.100 56.200 14.200 ;
        RECT 56.600 14.100 57.000 14.200 ;
        RECT 53.400 13.800 54.200 14.100 ;
        RECT 54.900 13.800 57.000 14.100 ;
        RECT 58.200 13.800 59.000 14.200 ;
        RECT 53.800 13.600 54.200 13.800 ;
        RECT 53.500 13.100 55.300 13.300 ;
        RECT 55.800 13.100 56.100 13.800 ;
        RECT 56.600 13.100 57.000 13.200 ;
        RECT 57.400 13.100 58.300 13.200 ;
        RECT 44.600 11.100 45.000 13.100 ;
        RECT 45.400 12.800 47.200 13.100 ;
        RECT 45.300 12.400 45.700 12.800 ;
        RECT 46.800 11.100 47.200 12.800 ;
        RECT 50.700 11.100 51.500 13.100 ;
        RECT 53.400 13.000 55.400 13.100 ;
        RECT 53.400 11.100 53.800 13.000 ;
        RECT 55.000 11.100 55.400 13.000 ;
        RECT 55.800 11.100 56.200 13.100 ;
        RECT 56.600 12.800 58.300 13.100 ;
        RECT 60.100 12.500 60.400 15.800 ;
        RECT 63.800 14.400 64.200 15.200 ;
        RECT 64.500 14.200 64.800 15.900 ;
        RECT 65.400 15.800 65.800 15.900 ;
        RECT 66.200 15.900 66.900 16.200 ;
        RECT 67.200 15.900 67.700 16.200 ;
        RECT 66.200 15.800 66.600 15.900 ;
        RECT 67.200 14.200 67.500 15.900 ;
        RECT 67.800 14.400 68.200 15.200 ;
        RECT 71.800 15.100 72.200 19.900 ;
        RECT 73.900 16.300 74.300 19.900 ;
        RECT 73.400 15.900 74.300 16.300 ;
        RECT 72.600 15.100 73.000 15.200 ;
        RECT 71.800 14.800 73.000 15.100 ;
        RECT 63.000 14.100 63.400 14.200 ;
        RECT 63.000 13.800 63.800 14.100 ;
        RECT 64.500 13.800 65.800 14.200 ;
        RECT 66.200 13.800 67.500 14.200 ;
        RECT 68.600 14.100 69.000 14.200 ;
        RECT 68.200 13.800 69.000 14.100 ;
        RECT 63.400 13.600 63.800 13.800 ;
        RECT 63.100 13.100 64.900 13.300 ;
        RECT 65.400 13.200 65.700 13.800 ;
        RECT 58.400 12.200 60.400 12.500 ;
        RECT 58.400 12.100 58.700 12.200 ;
        RECT 58.200 11.800 58.700 12.100 ;
        RECT 59.800 12.100 60.400 12.200 ;
        RECT 63.000 13.000 65.000 13.100 ;
        RECT 58.200 11.100 58.600 11.800 ;
        RECT 59.800 11.100 60.200 12.100 ;
        RECT 63.000 11.100 63.400 13.000 ;
        RECT 64.600 11.100 65.000 13.000 ;
        RECT 65.400 11.100 65.800 13.200 ;
        RECT 66.300 13.100 66.600 13.800 ;
        RECT 68.200 13.600 68.600 13.800 ;
        RECT 71.000 13.400 71.400 14.200 ;
        RECT 67.100 13.100 68.900 13.300 ;
        RECT 71.800 13.100 72.200 14.800 ;
        RECT 73.500 14.200 73.800 15.900 ;
        RECT 74.200 15.100 74.600 15.600 ;
        RECT 75.000 15.100 75.400 19.900 ;
        RECT 76.600 16.200 77.000 19.900 ;
        RECT 78.200 16.200 78.600 19.900 ;
        RECT 76.600 15.900 78.600 16.200 ;
        RECT 79.000 15.900 79.400 19.900 ;
        RECT 80.200 16.800 80.600 17.200 ;
        RECT 80.200 16.200 80.500 16.800 ;
        RECT 80.900 16.200 81.300 19.900 ;
        RECT 79.800 15.900 80.500 16.200 ;
        RECT 80.800 15.900 81.300 16.200 ;
        RECT 84.300 16.200 84.700 19.900 ;
        RECT 85.000 16.800 85.400 17.200 ;
        RECT 85.100 16.200 85.400 16.800 ;
        RECT 84.300 15.900 84.800 16.200 ;
        RECT 85.100 15.900 85.800 16.200 ;
        RECT 86.200 15.900 86.600 19.900 ;
        RECT 87.000 16.200 87.400 19.900 ;
        RECT 88.600 16.200 89.000 19.900 ;
        RECT 90.200 17.900 90.600 19.900 ;
        RECT 90.300 17.800 90.600 17.900 ;
        RECT 91.800 17.900 92.200 19.900 ;
        RECT 91.800 17.800 92.100 17.900 ;
        RECT 90.300 17.500 92.100 17.800 ;
        RECT 91.000 16.400 91.400 17.200 ;
        RECT 91.800 16.200 92.100 17.500 ;
        RECT 87.000 15.900 89.000 16.200 ;
        RECT 77.000 15.200 77.400 15.400 ;
        RECT 79.000 15.200 79.300 15.900 ;
        RECT 79.800 15.800 80.200 15.900 ;
        RECT 74.200 14.800 75.400 15.100 ;
        RECT 76.600 14.900 77.400 15.200 ;
        RECT 78.200 15.100 79.400 15.200 ;
        RECT 79.800 15.100 80.200 15.200 ;
        RECT 78.200 14.900 80.200 15.100 ;
        RECT 76.600 14.800 77.000 14.900 ;
        RECT 73.400 13.800 73.800 14.200 ;
        RECT 72.600 13.100 73.000 13.200 ;
        RECT 73.500 13.100 73.800 13.800 ;
        RECT 74.200 13.100 74.600 13.200 ;
        RECT 66.200 11.100 66.600 13.100 ;
        RECT 67.000 13.000 69.000 13.100 ;
        RECT 67.000 11.100 67.400 13.000 ;
        RECT 68.600 11.100 69.000 13.000 ;
        RECT 71.800 12.800 73.000 13.100 ;
        RECT 73.400 12.800 74.600 13.100 ;
        RECT 71.800 11.100 72.200 12.800 ;
        RECT 72.600 12.400 73.000 12.800 ;
        RECT 73.500 12.100 73.800 12.800 ;
        RECT 73.400 11.100 73.800 12.100 ;
        RECT 75.000 11.100 75.400 14.800 ;
        RECT 75.800 14.100 76.200 14.200 ;
        RECT 77.400 14.100 77.800 14.600 ;
        RECT 75.800 13.800 77.800 14.100 ;
        RECT 75.800 13.400 76.200 13.800 ;
        RECT 78.200 13.100 78.500 14.900 ;
        RECT 79.000 14.800 80.200 14.900 ;
        RECT 80.800 14.200 81.100 15.900 ;
        RECT 81.400 14.400 81.800 15.200 ;
        RECT 83.800 14.400 84.200 15.200 ;
        RECT 84.500 14.200 84.800 15.900 ;
        RECT 85.400 15.800 85.800 15.900 ;
        RECT 86.300 15.200 86.600 15.900 ;
        RECT 89.400 15.400 89.800 16.200 ;
        RECT 91.800 15.800 92.200 16.200 ;
        RECT 92.600 15.900 93.000 19.900 ;
        RECT 93.400 16.200 93.800 19.900 ;
        RECT 95.000 16.200 95.400 19.900 ;
        RECT 93.400 15.900 95.400 16.200 ;
        RECT 88.200 15.200 88.600 15.400 ;
        RECT 86.200 14.900 87.400 15.200 ;
        RECT 88.200 14.900 89.000 15.200 ;
        RECT 86.200 14.800 86.600 14.900 ;
        RECT 79.800 13.800 81.100 14.200 ;
        RECT 82.200 14.100 82.600 14.200 ;
        RECT 81.800 13.800 82.600 14.100 ;
        RECT 83.000 14.100 83.400 14.200 ;
        RECT 83.000 13.800 83.800 14.100 ;
        RECT 84.500 13.800 85.800 14.200 ;
        RECT 86.200 14.100 86.600 14.200 ;
        RECT 87.100 14.100 87.400 14.900 ;
        RECT 88.600 14.800 89.000 14.900 ;
        RECT 90.200 14.800 91.000 15.200 ;
        RECT 86.200 13.800 87.400 14.100 ;
        RECT 87.800 13.800 88.200 14.600 ;
        RECT 91.800 14.200 92.100 15.800 ;
        RECT 92.700 15.200 93.000 15.900 ;
        RECT 94.600 15.200 95.000 15.400 ;
        RECT 91.300 14.100 92.100 14.200 ;
        RECT 91.200 13.900 92.100 14.100 ;
        RECT 92.600 14.900 93.800 15.200 ;
        RECT 94.600 14.900 95.400 15.200 ;
        RECT 92.600 14.800 93.000 14.900 ;
        RECT 92.600 14.200 92.900 14.800 ;
        RECT 78.200 11.100 78.600 13.100 ;
        RECT 79.000 12.800 79.400 13.200 ;
        RECT 79.900 13.100 80.200 13.800 ;
        RECT 81.800 13.600 82.200 13.800 ;
        RECT 83.400 13.600 83.800 13.800 ;
        RECT 80.700 13.100 82.500 13.300 ;
        RECT 83.100 13.100 84.900 13.300 ;
        RECT 85.400 13.100 85.700 13.800 ;
        RECT 86.200 13.100 86.600 13.200 ;
        RECT 87.100 13.100 87.400 13.800 ;
        RECT 78.900 12.400 79.300 12.800 ;
        RECT 79.800 11.100 80.200 13.100 ;
        RECT 80.600 13.000 82.600 13.100 ;
        RECT 80.600 11.100 81.000 13.000 ;
        RECT 82.200 11.100 82.600 13.000 ;
        RECT 83.000 13.000 85.000 13.100 ;
        RECT 83.000 11.100 83.400 13.000 ;
        RECT 84.600 11.100 85.000 13.000 ;
        RECT 85.400 12.800 86.600 13.100 ;
        RECT 85.400 11.100 85.800 12.800 ;
        RECT 86.300 12.400 86.700 12.800 ;
        RECT 87.000 11.100 87.400 13.100 ;
        RECT 91.200 11.100 91.600 13.900 ;
        RECT 92.600 13.800 93.000 14.200 ;
        RECT 92.600 12.800 93.000 13.200 ;
        RECT 93.500 13.100 93.800 14.900 ;
        RECT 95.000 14.800 95.400 14.900 ;
        RECT 94.200 13.800 94.600 14.600 ;
        RECT 92.700 12.400 93.100 12.800 ;
        RECT 93.400 11.100 93.800 13.100 ;
        RECT 0.600 7.900 1.000 9.900 ;
        RECT 2.800 9.200 3.600 9.900 ;
        RECT 2.800 8.800 4.200 9.200 ;
        RECT 2.800 8.100 3.600 8.800 ;
        RECT 0.600 7.600 1.800 7.900 ;
        RECT 1.400 7.500 1.800 7.600 ;
        RECT 2.100 7.400 2.500 7.800 ;
        RECT 2.100 7.200 2.400 7.400 ;
        RECT 2.000 6.800 2.400 7.200 ;
        RECT 2.800 7.100 3.100 8.100 ;
        RECT 5.400 7.900 5.800 9.900 ;
        RECT 6.200 7.900 6.600 9.900 ;
        RECT 8.300 9.200 8.700 9.900 ;
        RECT 8.300 8.800 9.000 9.200 ;
        RECT 10.200 8.900 10.600 9.900 ;
        RECT 8.300 8.400 8.700 8.800 ;
        RECT 8.300 7.900 9.000 8.400 ;
        RECT 3.400 7.400 4.200 7.800 ;
        RECT 4.500 7.600 5.800 7.900 ;
        RECT 6.300 7.800 6.600 7.900 ;
        RECT 6.300 7.600 7.200 7.800 ;
        RECT 4.500 7.500 4.900 7.600 ;
        RECT 6.300 7.500 8.400 7.600 ;
        RECT 6.900 7.300 8.400 7.500 ;
        RECT 8.000 7.200 8.400 7.300 ;
        RECT 2.800 6.800 3.300 7.100 ;
        RECT 3.000 6.200 3.300 6.800 ;
        RECT 3.000 5.800 3.400 6.200 ;
        RECT 4.300 6.100 4.700 6.200 ;
        RECT 3.900 5.800 4.700 6.100 ;
        RECT 3.000 5.100 3.300 5.800 ;
        RECT 3.900 5.700 4.300 5.800 ;
        RECT 8.000 5.500 8.300 7.200 ;
        RECT 8.700 6.200 9.000 7.900 ;
        RECT 10.300 7.800 10.600 8.900 ;
        RECT 11.800 7.900 12.200 9.900 ;
        RECT 12.900 9.200 13.300 9.900 ;
        RECT 12.600 8.800 13.300 9.200 ;
        RECT 12.900 8.200 13.300 8.800 ;
        RECT 16.500 9.200 17.300 9.900 ;
        RECT 19.300 9.200 19.700 9.900 ;
        RECT 16.500 8.800 17.800 9.200 ;
        RECT 19.000 8.800 19.700 9.200 ;
        RECT 12.900 7.900 13.800 8.200 ;
        RECT 16.500 7.900 17.300 8.800 ;
        RECT 19.300 8.200 19.700 8.800 ;
        RECT 22.200 8.900 22.600 9.900 ;
        RECT 19.300 7.900 20.200 8.200 ;
        RECT 10.300 7.500 11.500 7.800 ;
        RECT 8.600 5.800 9.000 6.200 ;
        RECT 11.200 6.000 11.500 7.500 ;
        RECT 11.900 6.200 12.200 7.900 ;
        RECT 7.100 5.200 8.300 5.500 ;
        RECT 0.600 4.800 1.800 5.100 ;
        RECT 0.600 1.100 1.000 4.800 ;
        RECT 1.400 4.700 1.800 4.800 ;
        RECT 2.800 1.100 3.600 5.100 ;
        RECT 4.500 4.800 5.800 5.100 ;
        RECT 4.500 4.700 4.900 4.800 ;
        RECT 5.400 1.100 5.800 4.800 ;
        RECT 7.100 3.100 7.400 5.200 ;
        RECT 8.700 5.100 9.000 5.800 ;
        RECT 11.100 5.700 11.500 6.000 ;
        RECT 11.800 6.100 12.200 6.200 ;
        RECT 12.600 6.800 13.000 7.200 ;
        RECT 12.600 6.100 12.900 6.800 ;
        RECT 11.800 5.800 12.900 6.100 ;
        RECT 7.000 1.100 7.400 3.100 ;
        RECT 8.600 1.100 9.000 5.100 ;
        RECT 9.400 5.600 11.500 5.700 ;
        RECT 9.400 5.400 11.400 5.600 ;
        RECT 9.400 1.100 9.800 5.400 ;
        RECT 11.900 5.100 12.200 5.800 ;
        RECT 12.600 5.100 13.000 5.200 ;
        RECT 11.500 4.800 13.000 5.100 ;
        RECT 11.500 1.100 11.900 4.800 ;
        RECT 12.600 4.400 13.000 4.800 ;
        RECT 13.400 1.100 13.800 7.900 ;
        RECT 14.200 7.100 14.600 7.600 ;
        RECT 15.800 7.100 16.200 7.200 ;
        RECT 14.200 6.800 16.200 7.100 ;
        RECT 15.800 6.400 16.200 6.800 ;
        RECT 16.700 6.200 17.000 7.900 ;
        RECT 17.400 7.100 17.800 7.200 ;
        RECT 19.000 7.100 19.400 7.200 ;
        RECT 17.400 6.800 19.400 7.100 ;
        RECT 17.400 6.600 17.700 6.800 ;
        RECT 17.300 6.200 17.700 6.600 ;
        RECT 15.000 6.100 15.400 6.200 ;
        RECT 15.000 5.800 15.800 6.100 ;
        RECT 16.600 5.800 17.000 6.200 ;
        RECT 15.400 5.600 15.800 5.800 ;
        RECT 16.700 5.700 17.000 5.800 ;
        RECT 16.700 5.400 17.700 5.700 ;
        RECT 18.200 5.400 18.600 6.200 ;
        RECT 17.400 5.100 17.700 5.400 ;
        RECT 15.000 4.800 17.000 5.100 ;
        RECT 15.000 1.100 15.400 4.800 ;
        RECT 16.600 1.400 17.000 4.800 ;
        RECT 17.400 1.700 17.800 5.100 ;
        RECT 18.200 1.400 18.600 5.100 ;
        RECT 19.000 4.400 19.400 5.200 ;
        RECT 16.600 1.100 18.600 1.400 ;
        RECT 19.800 1.100 20.200 7.900 ;
        RECT 20.600 6.800 21.000 7.600 ;
        RECT 22.200 7.200 22.500 8.900 ;
        RECT 23.800 8.000 24.200 9.900 ;
        RECT 25.400 9.600 27.400 9.900 ;
        RECT 25.400 8.000 25.800 9.600 ;
        RECT 23.800 7.900 25.800 8.000 ;
        RECT 26.200 7.900 26.600 9.300 ;
        RECT 27.000 7.900 27.400 9.600 ;
        RECT 30.200 8.900 30.600 9.900 ;
        RECT 23.900 7.700 25.700 7.900 ;
        RECT 24.200 7.200 24.600 7.400 ;
        RECT 26.300 7.200 26.600 7.900 ;
        RECT 30.200 7.200 30.500 8.900 ;
        RECT 31.800 8.000 32.200 9.900 ;
        RECT 33.400 8.000 33.800 9.900 ;
        RECT 31.800 7.900 33.800 8.000 ;
        RECT 34.200 7.900 34.600 9.900 ;
        RECT 35.300 8.200 35.700 9.900 ;
        RECT 35.300 7.900 36.200 8.200 ;
        RECT 31.900 7.700 33.700 7.900 ;
        RECT 32.200 7.200 32.600 7.400 ;
        RECT 34.200 7.200 34.500 7.900 ;
        RECT 22.200 6.800 22.600 7.200 ;
        RECT 23.800 6.900 24.600 7.200 ;
        RECT 25.400 6.900 26.600 7.200 ;
        RECT 23.800 6.800 24.200 6.900 ;
        RECT 25.400 6.800 25.800 6.900 ;
        RECT 22.200 6.100 22.500 6.800 ;
        RECT 24.600 6.100 25.000 6.600 ;
        RECT 22.200 5.800 25.000 6.100 ;
        RECT 22.200 5.100 22.500 5.800 ;
        RECT 25.400 5.100 25.700 6.800 ;
        RECT 26.200 5.800 26.600 6.600 ;
        RECT 27.000 6.400 27.400 7.200 ;
        RECT 30.200 7.100 30.600 7.200 ;
        RECT 31.800 7.100 32.600 7.200 ;
        RECT 30.200 6.900 32.600 7.100 ;
        RECT 30.200 6.800 32.200 6.900 ;
        RECT 33.300 6.800 34.600 7.200 ;
        RECT 30.200 6.100 30.500 6.800 ;
        RECT 31.000 6.100 31.400 6.200 ;
        RECT 30.200 5.800 31.400 6.100 ;
        RECT 32.600 5.800 33.000 6.600 ;
        RECT 30.200 5.100 30.500 5.800 ;
        RECT 33.300 5.100 33.600 6.800 ;
        RECT 35.800 6.100 36.200 7.900 ;
        RECT 34.200 5.800 36.200 6.100 ;
        RECT 34.200 5.200 34.500 5.800 ;
        RECT 34.200 5.100 34.600 5.200 ;
        RECT 21.700 4.700 22.600 5.100 ;
        RECT 21.700 1.100 22.100 4.700 ;
        RECT 25.100 1.100 26.100 5.100 ;
        RECT 29.700 4.700 30.600 5.100 ;
        RECT 33.100 4.800 33.600 5.100 ;
        RECT 33.900 4.800 34.600 5.100 ;
        RECT 29.700 1.100 30.100 4.700 ;
        RECT 33.100 1.100 33.500 4.800 ;
        RECT 33.900 4.200 34.200 4.800 ;
        RECT 33.800 3.800 34.200 4.200 ;
        RECT 35.800 1.100 36.200 5.800 ;
        RECT 37.400 7.900 37.800 9.900 ;
        RECT 39.000 8.900 39.400 9.900 ;
        RECT 42.100 9.200 42.900 9.900 ;
        RECT 44.900 9.200 45.300 9.900 ;
        RECT 37.400 6.200 37.700 7.900 ;
        RECT 39.000 7.800 39.300 8.900 ;
        RECT 42.100 8.800 43.400 9.200 ;
        RECT 44.600 8.800 45.300 9.200 ;
        RECT 42.100 7.900 42.900 8.800 ;
        RECT 44.900 8.400 45.300 8.800 ;
        RECT 44.600 7.900 45.300 8.400 ;
        RECT 47.000 7.900 47.400 9.900 ;
        RECT 47.800 7.900 48.200 9.900 ;
        RECT 50.000 8.100 50.800 9.900 ;
        RECT 38.100 7.500 39.300 7.800 ;
        RECT 37.400 5.800 37.800 6.200 ;
        RECT 38.100 6.000 38.400 7.500 ;
        RECT 41.400 6.400 41.800 7.200 ;
        RECT 42.300 6.200 42.600 7.900 ;
        RECT 43.000 7.100 43.400 7.200 ;
        RECT 43.800 7.100 44.200 7.200 ;
        RECT 43.000 6.800 44.200 7.100 ;
        RECT 43.000 6.600 43.300 6.800 ;
        RECT 42.900 6.200 43.300 6.600 ;
        RECT 44.600 6.200 44.900 7.900 ;
        RECT 47.000 7.800 47.300 7.900 ;
        RECT 46.400 7.600 47.300 7.800 ;
        RECT 47.800 7.600 49.100 7.900 ;
        RECT 45.200 7.500 47.300 7.600 ;
        RECT 48.700 7.500 49.100 7.600 ;
        RECT 45.200 7.300 46.700 7.500 ;
        RECT 49.400 7.400 50.200 7.800 ;
        RECT 45.200 7.200 45.600 7.300 ;
        RECT 40.600 6.100 41.000 6.200 ;
        RECT 36.600 5.100 37.000 5.200 ;
        RECT 37.400 5.100 37.700 5.800 ;
        RECT 38.100 5.700 38.500 6.000 ;
        RECT 40.600 5.800 41.400 6.100 ;
        RECT 42.200 5.800 42.600 6.200 ;
        RECT 38.100 5.600 40.200 5.700 ;
        RECT 41.000 5.600 41.400 5.800 ;
        RECT 42.300 5.700 42.600 5.800 ;
        RECT 43.800 6.100 44.200 6.200 ;
        RECT 44.600 6.100 45.000 6.200 ;
        RECT 43.800 5.800 45.000 6.100 ;
        RECT 38.200 5.400 40.200 5.600 ;
        RECT 42.300 5.400 43.300 5.700 ;
        RECT 43.800 5.400 44.200 5.800 ;
        RECT 36.600 4.800 38.100 5.100 ;
        RECT 37.700 1.100 38.100 4.800 ;
        RECT 39.800 1.100 40.200 5.400 ;
        RECT 43.000 5.100 43.300 5.400 ;
        RECT 44.600 5.100 44.900 5.800 ;
        RECT 45.300 5.500 45.600 7.200 ;
        RECT 50.500 7.100 50.800 8.100 ;
        RECT 52.600 7.900 53.000 9.900 ;
        RECT 51.100 7.400 51.500 7.800 ;
        RECT 51.800 7.600 53.000 7.900 ;
        RECT 53.400 7.600 53.800 9.900 ;
        RECT 55.800 7.600 56.200 9.900 ;
        RECT 58.200 7.900 58.600 9.900 ;
        RECT 60.400 8.100 61.200 9.900 ;
        RECT 58.200 7.600 59.400 7.900 ;
        RECT 51.800 7.500 52.200 7.600 ;
        RECT 50.300 6.800 50.800 7.100 ;
        RECT 51.200 7.200 51.500 7.400 ;
        RECT 53.400 7.300 54.500 7.600 ;
        RECT 55.800 7.300 56.900 7.600 ;
        RECT 59.000 7.500 59.400 7.600 ;
        RECT 51.200 6.800 51.600 7.200 ;
        RECT 50.300 6.200 50.600 6.800 ;
        RECT 48.900 6.100 49.300 6.200 ;
        RECT 48.900 5.800 49.700 6.100 ;
        RECT 50.200 5.800 50.600 6.200 ;
        RECT 53.400 5.800 53.800 6.600 ;
        RECT 54.200 5.800 54.500 7.300 ;
        RECT 55.800 5.800 56.200 6.600 ;
        RECT 56.600 5.800 56.900 7.300 ;
        RECT 59.700 7.400 60.100 7.800 ;
        RECT 59.700 7.200 60.000 7.400 ;
        RECT 59.600 6.800 60.000 7.200 ;
        RECT 60.400 7.100 60.700 8.100 ;
        RECT 63.000 7.900 63.400 9.900 ;
        RECT 65.100 9.200 65.900 9.900 ;
        RECT 64.600 8.800 65.900 9.200 ;
        RECT 65.100 7.900 65.900 8.800 ;
        RECT 69.700 8.200 70.100 9.900 ;
        RECT 69.700 7.900 70.600 8.200 ;
        RECT 61.000 7.400 61.800 7.800 ;
        RECT 62.100 7.600 63.400 7.900 ;
        RECT 62.100 7.500 62.500 7.600 ;
        RECT 60.400 6.800 60.900 7.100 ;
        RECT 64.600 6.800 65.000 7.200 ;
        RECT 60.600 6.200 60.900 6.800 ;
        RECT 64.700 6.600 65.000 6.800 ;
        RECT 64.700 6.200 65.100 6.600 ;
        RECT 65.400 6.200 65.700 7.900 ;
        RECT 66.200 7.100 66.600 7.200 ;
        RECT 70.200 7.100 70.600 7.900 ;
        RECT 66.200 6.800 70.600 7.100 ;
        RECT 66.200 6.400 66.600 6.800 ;
        RECT 60.600 5.800 61.000 6.200 ;
        RECT 61.900 6.100 62.300 6.200 ;
        RECT 61.500 5.800 62.300 6.100 ;
        RECT 49.300 5.700 49.700 5.800 ;
        RECT 45.300 5.200 46.500 5.500 ;
        RECT 40.600 4.800 42.600 5.100 ;
        RECT 40.600 1.100 41.000 4.800 ;
        RECT 42.200 1.400 42.600 4.800 ;
        RECT 43.000 1.700 43.400 5.100 ;
        RECT 43.800 1.400 44.200 5.100 ;
        RECT 42.200 1.100 44.200 1.400 ;
        RECT 44.600 1.100 45.000 5.100 ;
        RECT 46.200 3.100 46.500 5.200 ;
        RECT 50.300 5.100 50.600 5.800 ;
        RECT 54.200 5.400 54.800 5.800 ;
        RECT 56.600 5.400 57.200 5.800 ;
        RECT 54.200 5.100 54.500 5.400 ;
        RECT 56.600 5.100 56.900 5.400 ;
        RECT 60.600 5.100 60.900 5.800 ;
        RECT 61.500 5.700 61.900 5.800 ;
        RECT 63.800 5.400 64.200 6.200 ;
        RECT 65.400 5.800 65.800 6.200 ;
        RECT 67.000 6.100 67.400 6.200 ;
        RECT 66.600 5.800 67.400 6.100 ;
        RECT 65.400 5.700 65.700 5.800 ;
        RECT 64.700 5.400 65.700 5.700 ;
        RECT 66.600 5.600 67.000 5.800 ;
        RECT 64.700 5.100 65.000 5.400 ;
        RECT 47.800 4.800 49.100 5.100 ;
        RECT 46.200 1.100 46.600 3.100 ;
        RECT 47.800 1.100 48.200 4.800 ;
        RECT 48.700 4.700 49.100 4.800 ;
        RECT 50.000 1.100 50.800 5.100 ;
        RECT 51.800 4.800 53.000 5.100 ;
        RECT 51.800 4.700 52.200 4.800 ;
        RECT 52.600 1.100 53.000 4.800 ;
        RECT 53.400 4.800 54.500 5.100 ;
        RECT 55.800 4.800 56.900 5.100 ;
        RECT 58.200 4.800 59.400 5.100 ;
        RECT 53.400 1.100 53.800 4.800 ;
        RECT 55.800 1.100 56.200 4.800 ;
        RECT 58.200 1.100 58.600 4.800 ;
        RECT 59.000 4.700 59.400 4.800 ;
        RECT 60.400 1.100 61.200 5.100 ;
        RECT 62.100 4.800 63.400 5.100 ;
        RECT 62.100 4.700 62.500 4.800 ;
        RECT 63.000 1.100 63.400 4.800 ;
        RECT 63.800 1.400 64.200 5.100 ;
        RECT 64.600 1.700 65.000 5.100 ;
        RECT 65.400 4.800 67.400 5.100 ;
        RECT 65.400 1.400 65.800 4.800 ;
        RECT 63.800 1.100 65.800 1.400 ;
        RECT 67.000 1.100 67.400 4.800 ;
        RECT 69.400 4.400 69.800 5.200 ;
        RECT 70.200 1.100 70.600 6.800 ;
        RECT 71.000 6.800 71.400 7.600 ;
        RECT 71.000 6.100 71.300 6.800 ;
        RECT 72.600 6.100 73.000 9.900 ;
        RECT 74.700 9.200 75.100 9.900 ;
        RECT 74.700 8.800 75.400 9.200 ;
        RECT 74.700 8.200 75.100 8.800 ;
        RECT 71.000 5.800 73.000 6.100 ;
        RECT 72.600 1.100 73.000 5.800 ;
        RECT 74.200 8.100 75.100 8.200 ;
        RECT 75.800 8.100 76.200 8.600 ;
        RECT 74.200 7.800 76.200 8.100 ;
        RECT 74.200 1.100 74.600 7.800 ;
        RECT 76.600 1.100 77.000 9.900 ;
        RECT 77.400 8.000 77.800 9.900 ;
        RECT 79.000 8.000 79.400 9.900 ;
        RECT 77.400 7.900 79.400 8.000 ;
        RECT 79.800 7.900 80.200 9.900 ;
        RECT 77.500 7.700 79.300 7.900 ;
        RECT 77.800 7.200 78.200 7.400 ;
        RECT 79.800 7.200 80.100 7.900 ;
        RECT 77.400 6.900 78.200 7.200 ;
        RECT 77.400 6.800 77.800 6.900 ;
        RECT 78.900 6.800 80.200 7.200 ;
        RECT 78.200 5.800 78.600 6.600 ;
        RECT 78.900 5.100 79.200 6.800 ;
        RECT 79.800 5.100 80.200 5.200 ;
        RECT 78.700 4.800 79.200 5.100 ;
        RECT 79.500 4.800 80.200 5.100 ;
        RECT 78.700 1.100 79.100 4.800 ;
        RECT 79.500 4.200 79.800 4.800 ;
        RECT 79.400 3.800 79.800 4.200 ;
        RECT 80.600 1.100 81.000 9.900 ;
        RECT 83.500 9.200 83.900 9.900 ;
        RECT 83.500 8.800 84.200 9.200 ;
        RECT 85.400 8.800 85.800 9.900 ;
        RECT 83.500 8.200 83.900 8.800 ;
        RECT 83.000 7.900 83.900 8.200 ;
        RECT 83.000 1.100 83.400 7.900 ;
        RECT 85.400 7.200 85.700 8.800 ;
        RECT 86.200 7.800 86.600 8.600 ;
        RECT 88.600 7.600 89.000 9.900 ;
        RECT 87.900 7.300 89.000 7.600 ;
        RECT 85.400 6.800 85.800 7.200 ;
        RECT 84.600 5.400 85.000 6.200 ;
        RECT 83.800 4.400 84.200 5.200 ;
        RECT 85.400 5.100 85.700 6.800 ;
        RECT 87.900 5.800 88.200 7.300 ;
        RECT 88.600 6.100 89.000 6.600 ;
        RECT 89.400 6.100 89.800 9.900 ;
        RECT 90.200 7.800 90.600 8.600 ;
        RECT 91.000 7.900 91.400 9.900 ;
        RECT 93.200 8.100 94.000 9.900 ;
        RECT 91.000 7.600 92.200 7.900 ;
        RECT 91.800 7.500 92.200 7.600 ;
        RECT 92.500 7.400 92.900 7.800 ;
        RECT 92.500 7.200 92.800 7.400 ;
        RECT 92.400 6.800 92.800 7.200 ;
        RECT 93.200 7.100 93.500 8.100 ;
        RECT 95.800 7.900 96.200 9.900 ;
        RECT 93.800 7.400 94.600 7.800 ;
        RECT 94.900 7.600 96.200 7.900 ;
        RECT 94.900 7.500 95.300 7.600 ;
        RECT 93.200 6.800 93.700 7.100 ;
        RECT 88.600 5.800 89.800 6.100 ;
        RECT 87.600 5.400 88.200 5.800 ;
        RECT 87.900 5.100 88.200 5.400 ;
        RECT 84.900 4.700 85.800 5.100 ;
        RECT 87.900 4.800 89.000 5.100 ;
        RECT 84.900 1.100 85.300 4.700 ;
        RECT 88.600 1.100 89.000 4.800 ;
        RECT 89.400 1.100 89.800 5.800 ;
        RECT 93.400 6.200 93.700 6.800 ;
        RECT 93.400 5.800 93.800 6.200 ;
        RECT 94.700 6.100 95.100 6.200 ;
        RECT 94.300 5.800 95.100 6.100 ;
        RECT 93.400 5.100 93.700 5.800 ;
        RECT 94.300 5.700 94.700 5.800 ;
        RECT 91.000 4.800 92.200 5.100 ;
        RECT 91.000 1.100 91.400 4.800 ;
        RECT 91.800 4.700 92.200 4.800 ;
        RECT 93.200 1.100 94.000 5.100 ;
        RECT 94.900 4.800 96.200 5.100 ;
        RECT 94.900 4.700 95.300 4.800 ;
        RECT 95.800 1.100 96.200 4.800 ;
      LAYER via1 ;
        RECT 3.800 72.800 4.200 73.200 ;
        RECT 13.400 76.800 13.800 77.200 ;
        RECT 11.800 74.800 12.200 75.200 ;
        RECT 7.000 71.800 7.400 72.200 ;
        RECT 10.200 71.800 10.600 72.200 ;
        RECT 16.600 71.800 17.000 72.200 ;
        RECT 25.400 74.800 25.800 75.200 ;
        RECT 21.400 71.800 21.800 72.200 ;
        RECT 31.000 71.800 31.400 72.200 ;
        RECT 38.200 76.800 38.600 77.200 ;
        RECT 39.800 76.800 40.200 77.200 ;
        RECT 35.800 73.800 36.200 74.200 ;
        RECT 35.000 71.800 35.400 72.200 ;
        RECT 44.600 74.800 45.000 75.200 ;
        RECT 39.000 71.800 39.400 72.200 ;
        RECT 44.600 72.800 45.000 73.200 ;
        RECT 45.400 71.800 45.800 72.200 ;
        RECT 47.000 71.800 47.400 72.200 ;
        RECT 53.400 73.800 53.800 74.200 ;
        RECT 55.000 73.800 55.400 74.200 ;
        RECT 52.600 72.800 53.000 73.200 ;
        RECT 71.800 76.800 72.200 77.200 ;
        RECT 61.400 74.800 61.800 75.200 ;
        RECT 70.200 75.800 70.600 76.200 ;
        RECT 67.000 74.800 67.400 75.200 ;
        RECT 67.800 73.800 68.200 74.200 ;
        RECT 75.800 76.800 76.200 77.200 ;
        RECT 74.200 74.800 74.600 75.200 ;
        RECT 59.800 71.800 60.200 72.200 ;
        RECT 76.600 74.800 77.000 75.200 ;
        RECT 78.200 74.800 78.600 75.200 ;
        RECT 74.200 72.800 74.600 73.200 ;
        RECT 81.400 72.800 81.800 73.200 ;
        RECT 90.200 74.800 90.600 75.200 ;
        RECT 92.600 74.800 93.000 75.200 ;
        RECT 96.600 74.800 97.000 75.200 ;
        RECT 4.600 68.800 5.000 69.200 ;
        RECT 5.400 67.800 5.800 68.200 ;
        RECT 4.600 66.800 5.000 67.200 ;
        RECT 3.800 65.800 4.200 66.200 ;
        RECT 7.000 64.800 7.400 65.200 ;
        RECT 9.400 65.800 9.800 66.200 ;
        RECT 13.400 65.800 13.800 66.200 ;
        RECT 15.000 64.800 15.400 65.200 ;
        RECT 17.400 64.800 17.800 65.200 ;
        RECT 15.800 62.800 16.200 63.200 ;
        RECT 22.200 65.800 22.600 66.200 ;
        RECT 23.800 65.800 24.200 66.200 ;
        RECT 26.200 65.800 26.600 66.200 ;
        RECT 30.200 65.800 30.600 66.200 ;
        RECT 29.400 64.800 29.800 65.200 ;
        RECT 32.600 65.800 33.000 66.200 ;
        RECT 35.000 65.800 35.400 66.200 ;
        RECT 42.200 65.800 42.600 66.200 ;
        RECT 21.400 61.800 21.800 62.200 ;
        RECT 26.200 61.800 26.600 62.200 ;
        RECT 32.600 61.800 33.000 62.200 ;
        RECT 35.000 61.800 35.400 62.200 ;
        RECT 37.400 61.800 37.800 62.200 ;
        RECT 47.000 66.800 47.400 67.200 ;
        RECT 53.400 66.800 53.800 67.200 ;
        RECT 44.600 65.800 45.000 66.200 ;
        RECT 47.800 65.800 48.200 66.200 ;
        RECT 43.800 62.800 44.200 63.200 ;
        RECT 50.200 64.800 50.600 65.200 ;
        RECT 55.000 66.800 55.400 67.200 ;
        RECT 63.000 66.800 63.400 67.200 ;
        RECT 55.800 65.800 56.200 66.200 ;
        RECT 53.400 61.800 53.800 62.200 ;
        RECT 59.000 65.800 59.400 66.200 ;
        RECT 65.400 65.800 65.800 66.200 ;
        RECT 58.200 61.800 58.600 62.200 ;
        RECT 65.400 63.800 65.800 64.200 ;
        RECT 71.000 65.800 71.400 66.200 ;
        RECT 70.200 62.800 70.600 63.200 ;
        RECT 68.600 61.800 69.000 62.200 ;
        RECT 90.200 68.800 90.600 69.200 ;
        RECT 74.200 64.800 74.600 65.200 ;
        RECT 77.400 64.800 77.800 65.200 ;
        RECT 79.800 65.800 80.200 66.200 ;
        RECT 82.200 65.800 82.600 66.200 ;
        RECT 84.600 65.800 85.000 66.200 ;
        RECT 87.800 66.800 88.200 67.200 ;
        RECT 88.600 65.800 89.000 66.200 ;
        RECT 92.600 68.800 93.000 69.200 ;
        RECT 91.000 66.800 91.400 67.200 ;
        RECT 91.800 65.800 92.200 66.200 ;
        RECT 84.600 62.800 85.000 63.200 ;
        RECT 96.600 65.800 97.000 66.200 ;
        RECT 94.200 64.800 94.600 65.200 ;
        RECT 95.000 61.800 95.400 62.200 ;
        RECT 5.400 58.800 5.800 59.200 ;
        RECT 4.600 56.800 5.000 57.200 ;
        RECT 10.200 54.800 10.600 55.200 ;
        RECT 14.200 55.800 14.600 56.200 ;
        RECT 11.800 54.800 12.200 55.200 ;
        RECT 8.600 51.800 9.000 52.200 ;
        RECT 10.200 51.800 10.600 52.200 ;
        RECT 25.400 58.800 25.800 59.200 ;
        RECT 22.200 56.800 22.600 57.200 ;
        RECT 18.200 54.800 18.600 55.200 ;
        RECT 16.600 51.800 17.000 52.200 ;
        RECT 26.200 53.800 26.600 54.200 ;
        RECT 34.200 57.800 34.600 58.200 ;
        RECT 48.600 58.800 49.000 59.200 ;
        RECT 41.400 54.800 41.800 55.200 ;
        RECT 46.200 54.800 46.600 55.200 ;
        RECT 41.400 53.800 41.800 54.200 ;
        RECT 43.800 52.800 44.200 53.200 ;
        RECT 47.000 53.800 47.400 54.200 ;
        RECT 44.600 51.800 45.000 52.200 ;
        RECT 47.800 52.800 48.200 53.200 ;
        RECT 53.400 54.800 53.800 55.200 ;
        RECT 56.600 54.800 57.000 55.200 ;
        RECT 51.000 53.800 51.400 54.200 ;
        RECT 58.200 53.800 58.600 54.200 ;
        RECT 61.400 54.800 61.800 55.200 ;
        RECT 73.400 58.800 73.800 59.200 ;
        RECT 74.200 56.800 74.600 57.200 ;
        RECT 50.200 52.800 50.600 53.200 ;
        RECT 63.800 53.800 64.200 54.200 ;
        RECT 59.800 52.800 60.200 53.200 ;
        RECT 59.000 51.800 59.400 52.200 ;
        RECT 61.400 52.800 61.800 53.200 ;
        RECT 69.400 54.800 69.800 55.200 ;
        RECT 65.400 52.800 65.800 53.200 ;
        RECT 66.200 52.800 66.600 53.200 ;
        RECT 67.000 51.800 67.400 52.200 ;
        RECT 72.600 55.800 73.000 56.200 ;
        RECT 87.800 58.800 88.200 59.200 ;
        RECT 82.200 54.800 82.600 55.200 ;
        RECT 87.800 54.800 88.200 55.200 ;
        RECT 71.800 52.800 72.200 53.200 ;
        RECT 75.800 52.800 76.200 53.200 ;
        RECT 83.000 53.800 83.400 54.200 ;
        RECT 85.400 52.800 85.800 53.200 ;
        RECT 88.600 53.800 89.000 54.200 ;
        RECT 91.000 58.800 91.400 59.200 ;
        RECT 92.600 54.800 93.000 55.200 ;
        RECT 95.800 54.800 96.200 55.200 ;
        RECT 96.600 53.800 97.000 54.200 ;
        RECT 3.800 48.800 4.200 49.200 ;
        RECT 7.000 48.800 7.400 49.200 ;
        RECT 10.200 48.800 10.600 49.200 ;
        RECT 3.800 44.800 4.200 45.200 ;
        RECT 7.000 44.800 7.400 45.200 ;
        RECT 15.800 45.800 16.200 46.200 ;
        RECT 13.400 41.800 13.800 42.200 ;
        RECT 27.000 44.800 27.400 45.200 ;
        RECT 30.200 44.800 30.600 45.200 ;
        RECT 32.600 45.800 33.000 46.200 ;
        RECT 35.800 45.800 36.200 46.200 ;
        RECT 33.400 41.800 33.800 42.200 ;
        RECT 43.800 46.800 44.200 47.200 ;
        RECT 49.400 46.800 49.800 47.200 ;
        RECT 39.000 45.800 39.400 46.200 ;
        RECT 42.200 45.800 42.600 46.200 ;
        RECT 38.200 44.800 38.600 45.200 ;
        RECT 47.800 45.800 48.200 46.200 ;
        RECT 50.200 48.800 50.600 49.200 ;
        RECT 55.800 48.800 56.200 49.200 ;
        RECT 52.600 46.800 53.000 47.200 ;
        RECT 56.600 46.800 57.000 47.200 ;
        RECT 71.000 48.800 71.400 49.200 ;
        RECT 63.800 46.800 64.200 47.200 ;
        RECT 70.200 46.800 70.600 47.200 ;
        RECT 50.200 41.800 50.600 42.200 ;
        RECT 59.000 44.800 59.400 45.200 ;
        RECT 67.800 45.800 68.200 46.200 ;
        RECT 67.000 44.800 67.400 45.200 ;
        RECT 81.400 46.800 81.800 47.200 ;
        RECT 79.000 45.800 79.400 46.200 ;
        RECT 90.200 48.800 90.600 49.200 ;
        RECT 83.800 46.800 84.200 47.200 ;
        RECT 85.400 46.800 85.800 47.200 ;
        RECT 83.000 45.800 83.400 46.200 ;
        RECT 76.600 43.800 77.000 44.200 ;
        RECT 75.000 42.800 75.400 43.200 ;
        RECT 79.800 44.800 80.200 45.200 ;
        RECT 85.400 45.800 85.800 46.200 ;
        RECT 97.400 48.800 97.800 49.200 ;
        RECT 91.000 46.800 91.400 47.200 ;
        RECT 89.400 45.800 89.800 46.200 ;
        RECT 1.400 34.800 1.800 35.200 ;
        RECT 8.600 34.800 9.000 35.200 ;
        RECT 3.000 31.800 3.400 32.200 ;
        RECT 15.000 32.800 15.400 33.200 ;
        RECT 11.800 31.800 12.200 32.200 ;
        RECT 13.400 31.800 13.800 32.200 ;
        RECT 29.400 34.800 29.800 35.200 ;
        RECT 23.800 33.800 24.200 34.200 ;
        RECT 19.800 31.800 20.200 32.200 ;
        RECT 43.800 38.800 44.200 39.200 ;
        RECT 47.000 36.800 47.400 37.200 ;
        RECT 52.600 36.800 53.000 37.200 ;
        RECT 33.400 33.800 33.800 34.200 ;
        RECT 38.200 34.800 38.600 35.200 ;
        RECT 32.600 31.800 33.000 32.200 ;
        RECT 35.800 31.800 36.200 32.200 ;
        RECT 41.400 32.800 41.800 33.200 ;
        RECT 42.200 32.800 42.600 33.200 ;
        RECT 49.400 32.800 49.800 33.200 ;
        RECT 55.800 34.800 56.200 35.200 ;
        RECT 55.000 33.800 55.400 34.200 ;
        RECT 56.600 33.800 57.000 34.200 ;
        RECT 62.200 34.800 62.600 35.200 ;
        RECT 66.200 34.800 66.600 35.200 ;
        RECT 63.000 33.800 63.400 34.200 ;
        RECT 67.000 33.800 67.400 34.200 ;
        RECT 63.800 32.800 64.200 33.200 ;
        RECT 76.600 34.800 77.000 35.200 ;
        RECT 85.400 38.800 85.800 39.200 ;
        RECT 87.000 38.800 87.400 39.200 ;
        RECT 63.000 31.800 63.400 32.200 ;
        RECT 74.200 31.800 74.600 32.200 ;
        RECT 79.000 32.800 79.400 33.200 ;
        RECT 82.200 34.800 82.600 35.200 ;
        RECT 86.200 34.800 86.600 35.200 ;
        RECT 83.000 33.800 83.400 34.200 ;
        RECT 86.200 33.800 86.600 34.200 ;
        RECT 95.000 35.800 95.400 36.200 ;
        RECT 89.400 34.800 89.800 35.200 ;
        RECT 90.200 34.800 90.600 35.200 ;
        RECT 87.800 33.800 88.200 34.200 ;
        RECT 15.800 28.800 16.200 29.200 ;
        RECT 11.800 26.800 12.200 27.200 ;
        RECT 3.000 24.800 3.400 25.200 ;
        RECT 16.600 26.800 17.000 27.200 ;
        RECT 19.000 26.800 19.400 27.200 ;
        RECT 15.000 25.800 15.400 26.200 ;
        RECT 7.000 21.800 7.400 22.200 ;
        RECT 37.400 28.800 37.800 29.200 ;
        RECT 23.000 22.800 23.400 23.200 ;
        RECT 29.400 25.800 29.800 26.200 ;
        RECT 27.000 24.800 27.400 25.200 ;
        RECT 33.400 25.800 33.800 26.200 ;
        RECT 41.400 25.800 41.800 26.200 ;
        RECT 43.800 25.800 44.200 26.200 ;
        RECT 47.800 26.800 48.200 27.200 ;
        RECT 44.600 24.800 45.000 25.200 ;
        RECT 50.200 25.800 50.600 26.200 ;
        RECT 58.200 28.800 58.600 29.200 ;
        RECT 61.400 28.800 61.800 29.200 ;
        RECT 55.000 26.800 55.400 27.200 ;
        RECT 57.400 26.800 57.800 27.200 ;
        RECT 49.400 22.800 49.800 23.200 ;
        RECT 55.800 25.800 56.200 26.200 ;
        RECT 60.600 26.800 61.000 27.200 ;
        RECT 65.400 24.800 65.800 25.200 ;
        RECT 73.400 24.800 73.800 25.200 ;
        RECT 76.600 26.800 77.000 27.200 ;
        RECT 79.000 26.800 79.400 27.200 ;
        RECT 82.200 26.800 82.600 27.200 ;
        RECT 89.400 24.800 89.800 25.200 ;
        RECT 87.800 23.800 88.200 24.200 ;
        RECT 91.800 25.800 92.200 26.200 ;
        RECT 92.600 21.800 93.000 22.200 ;
        RECT 9.400 16.800 9.800 17.200 ;
        RECT 11.000 16.800 11.400 17.200 ;
        RECT 3.800 14.800 4.200 15.200 ;
        RECT 12.600 15.800 13.000 16.200 ;
        RECT 11.800 14.800 12.200 15.200 ;
        RECT 15.000 16.800 15.400 17.200 ;
        RECT 3.000 13.800 3.400 14.200 ;
        RECT 4.600 13.800 5.000 14.200 ;
        RECT 5.400 12.800 5.800 13.200 ;
        RECT 13.400 13.800 13.800 14.200 ;
        RECT 23.000 14.800 23.400 15.200 ;
        RECT 19.800 12.800 20.200 13.200 ;
        RECT 23.800 13.800 24.200 14.200 ;
        RECT 28.600 13.800 29.000 14.200 ;
        RECT 33.400 18.800 33.800 19.200 ;
        RECT 31.000 15.800 31.400 16.200 ;
        RECT 47.000 16.800 47.400 17.200 ;
        RECT 26.200 11.800 26.600 12.200 ;
        RECT 37.400 12.800 37.800 13.200 ;
        RECT 36.600 11.800 37.000 12.200 ;
        RECT 40.600 11.800 41.000 12.200 ;
        RECT 48.600 15.800 49.000 16.200 ;
        RECT 61.400 17.800 61.800 18.200 ;
        RECT 47.800 14.800 48.200 15.200 ;
        RECT 54.200 14.800 54.600 15.200 ;
        RECT 56.600 13.800 57.000 14.200 ;
        RECT 63.800 14.800 64.200 15.200 ;
        RECT 67.800 14.800 68.200 15.200 ;
        RECT 75.000 18.800 75.400 19.200 ;
        RECT 72.600 14.800 73.000 15.200 ;
        RECT 65.400 12.800 65.800 13.200 ;
        RECT 68.600 13.800 69.000 14.200 ;
        RECT 71.000 13.800 71.400 14.200 ;
        RECT 66.200 11.800 66.600 12.200 ;
        RECT 74.200 12.800 74.600 13.200 ;
        RECT 79.800 14.800 80.200 15.200 ;
        RECT 81.400 14.800 81.800 15.200 ;
        RECT 83.800 14.800 84.200 15.200 ;
        RECT 90.200 18.800 90.600 19.200 ;
        RECT 91.000 16.800 91.400 17.200 ;
        RECT 89.400 15.800 89.800 16.200 ;
        RECT 82.200 13.800 82.600 14.200 ;
        RECT 79.800 11.800 80.200 12.200 ;
        RECT 3.800 8.800 4.200 9.200 ;
        RECT 8.600 8.800 9.000 9.200 ;
        RECT 3.800 7.400 4.200 7.800 ;
        RECT 17.400 8.800 17.800 9.200 ;
        RECT 15.800 6.800 16.200 7.200 ;
        RECT 19.000 6.800 19.400 7.200 ;
        RECT 18.200 5.800 18.600 6.200 ;
        RECT 19.000 4.800 19.400 5.200 ;
        RECT 27.000 6.800 27.400 7.200 ;
        RECT 33.400 6.800 33.800 7.200 ;
        RECT 31.000 5.800 31.400 6.200 ;
        RECT 34.200 4.800 34.600 5.200 ;
        RECT 43.000 8.800 43.400 9.200 ;
        RECT 50.200 8.800 50.600 9.200 ;
        RECT 41.400 6.800 41.800 7.200 ;
        RECT 43.800 6.800 44.200 7.200 ;
        RECT 60.600 8.800 61.000 9.200 ;
        RECT 61.400 7.400 61.800 7.800 ;
        RECT 63.800 5.800 64.200 6.200 ;
        RECT 67.000 5.800 67.400 6.200 ;
        RECT 69.400 4.800 69.800 5.200 ;
        RECT 75.000 8.800 75.400 9.200 ;
        RECT 76.600 8.800 77.000 9.200 ;
        RECT 72.600 5.800 73.000 6.200 ;
        RECT 79.000 6.800 79.400 7.200 ;
        RECT 83.800 8.800 84.200 9.200 ;
        RECT 80.600 5.800 81.000 6.200 ;
        RECT 79.800 4.800 80.200 5.200 ;
        RECT 84.600 5.800 85.000 6.200 ;
        RECT 83.800 4.800 84.200 5.200 ;
        RECT 93.400 8.800 93.800 9.200 ;
        RECT 94.200 7.400 94.600 7.800 ;
      LAYER metal2 ;
        RECT 39.800 77.800 40.200 78.200 ;
        RECT 71.000 77.800 71.400 78.200 ;
        RECT 39.800 77.200 40.100 77.800 ;
        RECT 13.400 76.800 13.800 77.200 ;
        RECT 37.400 76.800 37.800 77.200 ;
        RECT 38.200 77.100 38.600 77.200 ;
        RECT 39.000 77.100 39.400 77.200 ;
        RECT 38.200 76.800 39.400 77.100 ;
        RECT 39.800 76.800 40.200 77.200 ;
        RECT 13.400 76.200 13.700 76.800 ;
        RECT 11.800 75.800 12.200 76.200 ;
        RECT 13.400 75.800 13.800 76.200 ;
        RECT 16.600 76.100 17.000 76.200 ;
        RECT 17.400 76.100 17.800 76.200 ;
        RECT 16.600 75.800 17.800 76.100 ;
        RECT 19.000 75.800 19.400 76.200 ;
        RECT 25.400 75.800 25.800 76.200 ;
        RECT 26.200 76.100 26.600 76.200 ;
        RECT 27.000 76.100 27.400 76.200 ;
        RECT 26.200 75.800 27.400 76.100 ;
        RECT 11.800 75.200 12.100 75.800 ;
        RECT 16.600 75.200 16.900 75.800 ;
        RECT 19.000 75.200 19.300 75.800 ;
        RECT 25.400 75.200 25.700 75.800 ;
        RECT 37.400 75.200 37.700 76.800 ;
        RECT 71.000 76.200 71.300 77.800 ;
        RECT 71.800 77.100 72.200 77.200 ;
        RECT 72.600 77.100 73.000 77.200 ;
        RECT 71.800 76.800 73.000 77.100 ;
        RECT 75.800 77.100 76.200 77.200 ;
        RECT 76.600 77.100 77.000 77.200 ;
        RECT 75.800 76.800 77.000 77.100 ;
        RECT 64.600 75.800 65.000 76.200 ;
        RECT 65.400 75.800 65.800 76.200 ;
        RECT 70.200 75.800 70.600 76.200 ;
        RECT 71.000 75.800 71.400 76.200 ;
        RECT 64.600 75.200 64.900 75.800 ;
        RECT 11.800 74.800 12.200 75.200 ;
        RECT 16.600 74.800 17.000 75.200 ;
        RECT 19.000 74.800 19.400 75.200 ;
        RECT 25.400 74.800 25.800 75.200 ;
        RECT 37.400 74.800 37.800 75.200 ;
        RECT 44.600 74.800 45.000 75.200 ;
        RECT 51.000 74.800 51.400 75.200 ;
        RECT 61.400 74.800 61.800 75.200 ;
        RECT 64.600 74.800 65.000 75.200 ;
        RECT 35.800 73.800 36.200 74.200 ;
        RECT 35.800 73.200 36.100 73.800 ;
        RECT 37.400 73.200 37.700 74.800 ;
        RECT 44.600 73.200 44.900 74.800 ;
        RECT 3.800 72.800 4.200 73.200 ;
        RECT 23.800 72.800 24.200 73.200 ;
        RECT 28.600 72.800 29.000 73.200 ;
        RECT 35.800 72.800 36.200 73.200 ;
        RECT 37.400 72.800 37.800 73.200 ;
        RECT 44.600 72.800 45.000 73.200 ;
        RECT 49.400 73.100 49.800 73.200 ;
        RECT 50.200 73.100 50.600 73.200 ;
        RECT 49.400 72.800 50.600 73.100 ;
        RECT 3.800 69.100 4.100 72.800 ;
        RECT 7.000 71.800 7.400 72.200 ;
        RECT 10.200 71.800 10.600 72.200 ;
        RECT 15.800 72.100 16.200 72.200 ;
        RECT 16.600 72.100 17.000 72.200 ;
        RECT 15.800 71.800 17.000 72.100 ;
        RECT 21.400 71.800 21.800 72.200 ;
        RECT 7.000 69.200 7.300 71.800 ;
        RECT 4.600 69.100 5.000 69.200 ;
        RECT 5.400 69.100 5.800 69.200 ;
        RECT 3.800 68.800 5.800 69.100 ;
        RECT 7.000 68.800 7.400 69.200 ;
        RECT 10.200 68.200 10.500 71.800 ;
        RECT 21.400 71.200 21.700 71.800 ;
        RECT 21.400 70.800 21.800 71.200 ;
        RECT 22.200 69.800 22.600 70.200 ;
        RECT 4.600 67.800 5.000 68.200 ;
        RECT 5.400 67.800 5.800 68.200 ;
        RECT 10.200 67.800 10.600 68.200 ;
        RECT 11.000 67.800 11.400 68.200 ;
        RECT 19.000 68.100 19.400 68.200 ;
        RECT 19.800 68.100 20.200 68.200 ;
        RECT 19.000 67.800 20.200 68.100 ;
        RECT 4.600 67.200 4.900 67.800 ;
        RECT 4.600 66.800 5.000 67.200 ;
        RECT 3.800 65.800 4.200 66.200 ;
        RECT 3.800 60.200 4.100 65.800 ;
        RECT 3.800 59.800 4.200 60.200 ;
        RECT 5.400 59.200 5.700 67.800 ;
        RECT 8.600 65.800 9.000 66.200 ;
        RECT 9.400 65.800 9.800 66.200 ;
        RECT 8.600 65.200 8.900 65.800 ;
        RECT 7.000 64.800 7.400 65.200 ;
        RECT 8.600 64.800 9.000 65.200 ;
        RECT 7.000 64.200 7.300 64.800 ;
        RECT 7.000 63.800 7.400 64.200 ;
        RECT 5.400 58.800 5.800 59.200 ;
        RECT 4.600 56.800 5.000 57.200 ;
        RECT 2.200 55.800 2.600 56.200 ;
        RECT 0.600 45.800 1.000 46.200 ;
        RECT 0.600 34.200 0.900 45.800 ;
        RECT 2.200 43.200 2.500 55.800 ;
        RECT 3.800 54.800 4.200 55.200 ;
        RECT 3.800 49.200 4.100 54.800 ;
        RECT 4.600 53.200 4.900 56.800 ;
        RECT 9.400 54.200 9.700 65.800 ;
        RECT 10.200 54.800 10.600 55.200 ;
        RECT 9.400 53.800 9.800 54.200 ;
        RECT 4.600 52.800 5.000 53.200 ;
        RECT 7.000 52.800 7.400 53.200 ;
        RECT 7.000 49.200 7.300 52.800 ;
        RECT 8.600 51.800 9.000 52.200 ;
        RECT 8.600 51.200 8.900 51.800 ;
        RECT 8.600 50.800 9.000 51.200 ;
        RECT 9.400 49.200 9.700 53.800 ;
        RECT 10.200 53.200 10.500 54.800 ;
        RECT 11.000 53.200 11.300 67.800 ;
        RECT 11.800 67.100 12.200 67.200 ;
        RECT 12.600 67.100 13.000 67.200 ;
        RECT 11.800 66.800 13.000 67.100 ;
        RECT 16.600 66.800 17.000 67.200 ;
        RECT 17.400 66.800 17.800 67.200 ;
        RECT 12.600 66.100 13.000 66.200 ;
        RECT 13.400 66.100 13.800 66.200 ;
        RECT 12.600 65.800 13.800 66.100 ;
        RECT 14.200 65.800 14.600 66.200 ;
        RECT 14.200 65.200 14.500 65.800 ;
        RECT 14.200 64.800 14.600 65.200 ;
        RECT 15.000 64.800 15.400 65.200 ;
        RECT 15.000 64.200 15.300 64.800 ;
        RECT 12.600 63.800 13.000 64.200 ;
        RECT 15.000 63.800 15.400 64.200 ;
        RECT 15.800 63.800 16.200 64.200 ;
        RECT 12.600 63.200 12.900 63.800 ;
        RECT 15.800 63.200 16.100 63.800 ;
        RECT 12.600 62.800 13.000 63.200 ;
        RECT 15.800 62.800 16.200 63.200 ;
        RECT 11.800 57.800 12.200 58.200 ;
        RECT 11.800 55.200 12.100 57.800 ;
        RECT 14.200 56.800 14.600 57.200 ;
        RECT 14.200 56.200 14.500 56.800 ;
        RECT 14.200 55.800 14.600 56.200 ;
        RECT 11.800 54.800 12.200 55.200 ;
        RECT 16.600 53.200 16.900 66.800 ;
        RECT 17.400 66.200 17.700 66.800 ;
        RECT 22.200 66.200 22.500 69.800 ;
        RECT 23.800 69.200 24.100 72.800 ;
        RECT 26.200 71.800 26.600 72.200 ;
        RECT 23.800 68.800 24.200 69.200 ;
        RECT 24.600 68.800 25.000 69.200 ;
        RECT 23.800 68.200 24.100 68.800 ;
        RECT 24.600 68.200 24.900 68.800 ;
        RECT 23.800 67.800 24.200 68.200 ;
        RECT 24.600 67.800 25.000 68.200 ;
        RECT 26.200 67.200 26.500 71.800 ;
        RECT 28.600 68.200 28.900 72.800 ;
        RECT 51.000 72.200 51.300 74.800 ;
        RECT 53.400 74.100 53.800 74.200 ;
        RECT 54.200 74.100 54.600 74.200 ;
        RECT 53.400 73.800 54.600 74.100 ;
        RECT 55.000 73.800 55.400 74.200 ;
        RECT 52.600 73.100 53.000 73.200 ;
        RECT 53.400 73.100 53.800 73.200 ;
        RECT 52.600 72.800 53.800 73.100 ;
        RECT 30.200 71.800 30.600 72.200 ;
        RECT 31.000 71.800 31.400 72.200 ;
        RECT 35.000 71.800 35.400 72.200 ;
        RECT 35.800 71.800 36.200 72.200 ;
        RECT 39.000 71.800 39.400 72.200 ;
        RECT 45.400 71.800 45.800 72.200 ;
        RECT 47.000 71.800 47.400 72.200 ;
        RECT 51.000 71.800 51.400 72.200 ;
        RECT 30.200 68.200 30.500 71.800 ;
        RECT 31.000 70.200 31.300 71.800 ;
        RECT 31.000 69.800 31.400 70.200 ;
        RECT 35.000 68.200 35.300 71.800 ;
        RECT 35.800 68.200 36.100 71.800 ;
        RECT 37.400 69.800 37.800 70.200 ;
        RECT 28.600 67.800 29.000 68.200 ;
        RECT 30.200 67.800 30.600 68.200 ;
        RECT 32.600 67.800 33.000 68.200 ;
        RECT 35.000 67.800 35.400 68.200 ;
        RECT 35.800 67.800 36.200 68.200 ;
        RECT 32.600 67.200 32.900 67.800 ;
        RECT 26.200 66.800 26.600 67.200 ;
        RECT 30.200 66.800 30.600 67.200 ;
        RECT 32.600 66.800 33.000 67.200 ;
        RECT 26.200 66.200 26.500 66.800 ;
        RECT 30.200 66.200 30.500 66.800 ;
        RECT 32.600 66.200 32.900 66.800 ;
        RECT 35.000 66.200 35.300 67.800 ;
        RECT 37.400 66.200 37.700 69.800 ;
        RECT 39.000 69.200 39.300 71.800 ;
        RECT 39.000 68.800 39.400 69.200 ;
        RECT 39.000 68.100 39.400 68.200 ;
        RECT 39.800 68.100 40.200 68.200 ;
        RECT 39.000 67.800 40.200 68.100 ;
        RECT 42.200 67.800 42.600 68.200 ;
        RECT 42.200 66.200 42.500 67.800 ;
        RECT 45.400 67.200 45.700 71.800 ;
        RECT 47.000 68.100 47.300 71.800 ;
        RECT 50.200 70.800 50.600 71.200 ;
        RECT 47.800 68.100 48.200 68.200 ;
        RECT 47.000 67.800 48.200 68.100 ;
        RECT 43.000 66.800 43.400 67.200 ;
        RECT 45.400 66.800 45.800 67.200 ;
        RECT 47.000 66.800 47.400 67.200 ;
        RECT 17.400 65.800 17.800 66.200 ;
        RECT 22.200 65.800 22.600 66.200 ;
        RECT 23.800 66.100 24.200 66.200 ;
        RECT 24.600 66.100 25.000 66.200 ;
        RECT 23.800 65.800 25.000 66.100 ;
        RECT 26.200 65.800 26.600 66.200 ;
        RECT 30.200 65.800 30.600 66.200 ;
        RECT 32.600 65.800 33.000 66.200 ;
        RECT 35.000 65.800 35.400 66.200 ;
        RECT 37.400 65.800 37.800 66.200 ;
        RECT 42.200 65.800 42.600 66.200 ;
        RECT 17.400 64.800 17.800 65.200 ;
        RECT 22.200 64.800 22.600 65.200 ;
        RECT 29.400 64.800 29.800 65.200 ;
        RECT 17.400 62.200 17.700 64.800 ;
        RECT 22.200 64.200 22.500 64.800 ;
        RECT 22.200 63.800 22.600 64.200 ;
        RECT 21.400 62.800 21.800 63.200 ;
        RECT 21.400 62.200 21.700 62.800 ;
        RECT 17.400 61.800 17.800 62.200 ;
        RECT 21.400 61.800 21.800 62.200 ;
        RECT 26.200 61.800 26.600 62.200 ;
        RECT 21.400 61.200 21.700 61.800 ;
        RECT 21.400 60.800 21.800 61.200 ;
        RECT 25.400 59.800 25.800 60.200 ;
        RECT 25.400 59.200 25.700 59.800 ;
        RECT 25.400 58.800 25.800 59.200 ;
        RECT 26.200 59.100 26.500 61.800 ;
        RECT 26.200 58.800 27.300 59.100 ;
        RECT 22.200 56.800 22.600 57.200 ;
        RECT 22.200 56.200 22.500 56.800 ;
        RECT 19.800 56.100 20.200 56.200 ;
        RECT 19.800 55.800 20.900 56.100 ;
        RECT 22.200 55.800 22.600 56.200 ;
        RECT 18.200 54.800 18.600 55.200 ;
        RECT 17.400 53.800 17.800 54.200 ;
        RECT 17.400 53.200 17.700 53.800 ;
        RECT 10.200 52.800 10.600 53.200 ;
        RECT 11.000 52.800 11.400 53.200 ;
        RECT 11.800 52.800 12.200 53.200 ;
        RECT 13.400 52.800 13.800 53.200 ;
        RECT 16.600 52.800 17.000 53.200 ;
        RECT 17.400 52.800 17.800 53.200 ;
        RECT 10.200 51.800 10.600 52.200 ;
        RECT 10.200 51.200 10.500 51.800 ;
        RECT 10.200 50.800 10.600 51.200 ;
        RECT 3.800 48.800 4.200 49.200 ;
        RECT 7.000 48.800 7.400 49.200 ;
        RECT 9.400 48.800 9.800 49.200 ;
        RECT 10.200 49.100 10.600 49.200 ;
        RECT 11.000 49.100 11.400 49.200 ;
        RECT 10.200 48.800 11.400 49.100 ;
        RECT 11.800 48.200 12.100 52.800 ;
        RECT 13.400 49.200 13.700 52.800 ;
        RECT 15.800 51.800 16.200 52.200 ;
        RECT 16.600 51.800 17.000 52.200 ;
        RECT 15.800 49.200 16.100 51.800 ;
        RECT 16.600 51.200 16.900 51.800 ;
        RECT 16.600 50.800 17.000 51.200 ;
        RECT 13.400 48.800 13.800 49.200 ;
        RECT 15.800 48.800 16.200 49.200 ;
        RECT 13.400 48.200 13.700 48.800 ;
        RECT 11.000 48.100 11.400 48.200 ;
        RECT 11.800 48.100 12.200 48.200 ;
        RECT 11.000 47.800 12.200 48.100 ;
        RECT 13.400 47.800 13.800 48.200 ;
        RECT 15.800 46.200 16.100 48.800 ;
        RECT 18.200 48.200 18.500 54.800 ;
        RECT 20.600 52.200 20.900 55.800 ;
        RECT 21.400 54.800 21.800 55.200 ;
        RECT 21.400 54.200 21.700 54.800 ;
        RECT 21.400 53.800 21.800 54.200 ;
        RECT 24.600 53.800 25.000 54.200 ;
        RECT 26.200 53.800 26.600 54.200 ;
        RECT 20.600 51.800 21.000 52.200 ;
        RECT 18.200 47.800 18.600 48.200 ;
        RECT 19.800 47.800 20.200 48.200 ;
        RECT 19.800 47.200 20.100 47.800 ;
        RECT 19.800 46.800 20.200 47.200 ;
        RECT 20.600 46.200 20.900 51.800 ;
        RECT 24.600 49.200 24.900 53.800 ;
        RECT 26.200 50.200 26.500 53.800 ;
        RECT 26.200 49.800 26.600 50.200 ;
        RECT 27.000 49.200 27.300 58.800 ;
        RECT 28.600 54.800 29.000 55.200 ;
        RECT 28.600 49.200 28.900 54.800 ;
        RECT 23.800 48.800 24.200 49.200 ;
        RECT 24.600 48.800 25.000 49.200 ;
        RECT 27.000 48.800 27.400 49.200 ;
        RECT 28.600 48.800 29.000 49.200 ;
        RECT 23.800 46.200 24.100 48.800 ;
        RECT 4.600 45.800 5.000 46.200 ;
        RECT 15.800 45.800 16.200 46.200 ;
        RECT 20.600 45.800 21.000 46.200 ;
        RECT 23.800 45.800 24.200 46.200 ;
        RECT 3.800 45.100 4.200 45.200 ;
        RECT 4.600 45.100 4.900 45.800 ;
        RECT 3.800 44.800 4.900 45.100 ;
        RECT 2.200 42.800 2.600 43.200 ;
        RECT 1.400 40.800 1.800 41.200 ;
        RECT 1.400 35.200 1.700 40.800 ;
        RECT 3.000 36.100 3.400 36.200 ;
        RECT 3.800 36.100 4.200 36.200 ;
        RECT 3.000 35.800 4.200 36.100 ;
        RECT 1.400 34.800 1.800 35.200 ;
        RECT 3.800 34.800 4.200 35.200 ;
        RECT 3.800 34.200 4.100 34.800 ;
        RECT 4.600 34.200 4.900 44.800 ;
        RECT 7.000 44.800 7.400 45.200 ;
        RECT 23.800 44.800 24.200 45.200 ;
        RECT 27.000 45.100 27.400 45.200 ;
        RECT 27.800 45.100 28.200 45.200 ;
        RECT 27.000 44.800 28.200 45.100 ;
        RECT 7.000 44.200 7.300 44.800 ;
        RECT 23.800 44.200 24.100 44.800 ;
        RECT 7.000 43.800 7.400 44.200 ;
        RECT 16.600 44.100 17.000 44.200 ;
        RECT 17.400 44.100 17.800 44.200 ;
        RECT 16.600 43.800 17.800 44.100 ;
        RECT 23.800 43.800 24.200 44.200 ;
        RECT 24.600 44.100 25.000 44.200 ;
        RECT 25.400 44.100 25.800 44.200 ;
        RECT 24.600 43.800 25.800 44.100 ;
        RECT 29.400 43.200 29.700 64.800 ;
        RECT 37.400 64.100 37.800 64.200 ;
        RECT 38.200 64.100 38.600 64.200 ;
        RECT 37.400 63.800 38.600 64.100 ;
        RECT 43.000 63.200 43.300 66.800 ;
        RECT 43.800 66.100 44.200 66.200 ;
        RECT 44.600 66.100 45.000 66.200 ;
        RECT 43.800 65.800 45.000 66.100 ;
        RECT 46.200 65.800 46.600 66.200 ;
        RECT 46.200 65.200 46.500 65.800 ;
        RECT 46.200 64.800 46.600 65.200 ;
        RECT 43.000 62.800 43.400 63.200 ;
        RECT 43.800 63.100 44.200 63.200 ;
        RECT 44.600 63.100 45.000 63.200 ;
        RECT 43.800 62.800 45.000 63.100 ;
        RECT 32.600 62.100 33.000 62.200 ;
        RECT 33.400 62.100 33.800 62.200 ;
        RECT 32.600 61.800 33.800 62.100 ;
        RECT 35.000 61.800 35.400 62.200 ;
        RECT 37.400 62.100 37.800 62.200 ;
        RECT 37.400 61.800 38.500 62.100 ;
        RECT 35.000 61.200 35.300 61.800 ;
        RECT 35.000 60.800 35.400 61.200 ;
        RECT 35.000 59.200 35.300 60.800 ;
        RECT 35.000 58.800 35.400 59.200 ;
        RECT 34.200 57.800 34.600 58.200 ;
        RECT 34.200 57.200 34.500 57.800 ;
        RECT 34.200 56.800 34.600 57.200 ;
        RECT 37.400 56.800 37.800 57.200 ;
        RECT 31.000 56.100 31.400 56.200 ;
        RECT 31.800 56.100 32.200 56.200 ;
        RECT 31.000 55.800 32.200 56.100 ;
        RECT 35.000 55.800 35.400 56.200 ;
        RECT 31.000 51.200 31.300 55.800 ;
        RECT 35.000 55.200 35.300 55.800 ;
        RECT 35.000 55.100 35.400 55.200 ;
        RECT 35.000 54.800 36.100 55.100 ;
        RECT 31.000 50.800 31.400 51.200 ;
        RECT 35.800 48.200 36.100 54.800 ;
        RECT 36.600 54.800 37.000 55.200 ;
        RECT 36.600 54.200 36.900 54.800 ;
        RECT 37.400 54.200 37.700 56.800 ;
        RECT 36.600 53.800 37.000 54.200 ;
        RECT 37.400 53.800 37.800 54.200 ;
        RECT 38.200 51.200 38.500 61.800 ;
        RECT 39.800 61.800 40.200 62.200 ;
        RECT 41.400 61.800 41.800 62.200 ;
        RECT 39.800 56.200 40.100 61.800 ;
        RECT 39.000 55.800 39.400 56.200 ;
        RECT 39.800 55.800 40.200 56.200 ;
        RECT 39.000 52.200 39.300 55.800 ;
        RECT 39.000 51.800 39.400 52.200 ;
        RECT 38.200 50.800 38.600 51.200 ;
        RECT 37.400 49.800 37.800 50.200 ;
        RECT 37.400 49.200 37.700 49.800 ;
        RECT 37.400 48.800 37.800 49.200 ;
        RECT 35.800 47.800 36.200 48.200 ;
        RECT 31.800 46.800 32.200 47.200 ;
        RECT 31.800 45.200 32.100 46.800 ;
        RECT 35.800 46.200 36.100 47.800 ;
        RECT 36.600 46.800 37.000 47.200 ;
        RECT 32.600 45.800 33.000 46.200 ;
        RECT 35.800 45.800 36.200 46.200 ;
        RECT 30.200 44.800 30.600 45.200 ;
        RECT 31.800 44.800 32.200 45.200 ;
        RECT 30.200 44.200 30.500 44.800 ;
        RECT 32.600 44.200 32.900 45.800 ;
        RECT 30.200 43.800 30.600 44.200 ;
        RECT 32.600 43.800 33.000 44.200 ;
        RECT 29.400 42.800 29.800 43.200 ;
        RECT 29.400 42.200 29.700 42.800 ;
        RECT 13.400 41.800 13.800 42.200 ;
        RECT 20.600 41.800 21.000 42.200 ;
        RECT 29.400 41.800 29.800 42.200 ;
        RECT 33.400 41.800 33.800 42.200 ;
        RECT 7.000 40.800 7.400 41.200 ;
        RECT 5.400 35.800 5.800 36.200 ;
        RECT 5.400 35.200 5.700 35.800 ;
        RECT 7.000 35.200 7.300 40.800 ;
        RECT 8.600 38.800 9.000 39.200 ;
        RECT 8.600 35.200 8.900 38.800 ;
        RECT 11.800 36.800 12.200 37.200 ;
        RECT 11.800 36.200 12.100 36.800 ;
        RECT 9.400 35.800 9.800 36.200 ;
        RECT 11.800 35.800 12.200 36.200 ;
        RECT 5.400 34.800 5.800 35.200 ;
        RECT 7.000 34.800 7.400 35.200 ;
        RECT 7.800 35.100 8.200 35.200 ;
        RECT 8.600 35.100 9.000 35.200 ;
        RECT 7.800 34.800 9.000 35.100 ;
        RECT 9.400 34.200 9.700 35.800 ;
        RECT 13.400 35.200 13.700 41.800 ;
        RECT 20.600 38.200 20.900 41.800 ;
        RECT 24.600 38.800 25.000 39.200 ;
        RECT 20.600 37.800 21.000 38.200 ;
        RECT 19.000 36.800 19.400 37.200 ;
        RECT 14.200 36.100 14.600 36.200 ;
        RECT 14.200 35.800 15.300 36.100 ;
        RECT 14.200 35.200 14.500 35.800 ;
        RECT 13.400 34.800 13.800 35.200 ;
        RECT 14.200 34.800 14.600 35.200 ;
        RECT 0.600 33.800 1.000 34.200 ;
        RECT 3.800 33.800 4.200 34.200 ;
        RECT 4.600 33.800 5.000 34.200 ;
        RECT 6.200 33.800 6.600 34.200 ;
        RECT 9.400 33.800 9.800 34.200 ;
        RECT 0.600 33.200 0.900 33.800 ;
        RECT 0.600 32.800 1.000 33.200 ;
        RECT 3.000 31.800 3.400 32.200 ;
        RECT 3.000 26.100 3.300 31.800 ;
        RECT 6.200 31.200 6.500 33.800 ;
        RECT 9.400 33.200 9.700 33.800 ;
        RECT 15.000 33.200 15.300 35.800 ;
        RECT 16.600 35.800 17.000 36.200 ;
        RECT 9.400 32.800 9.800 33.200 ;
        RECT 15.000 32.800 15.400 33.200 ;
        RECT 11.800 31.800 12.200 32.200 ;
        RECT 13.400 31.800 13.800 32.200 ;
        RECT 6.200 30.800 6.600 31.200 ;
        RECT 6.200 29.800 6.600 30.200 ;
        RECT 4.600 27.100 5.000 27.200 ;
        RECT 5.400 27.100 5.800 27.200 ;
        RECT 4.600 26.800 5.800 27.100 ;
        RECT 6.200 26.200 6.500 29.800 ;
        RECT 10.200 27.800 10.600 28.200 ;
        RECT 8.600 27.100 9.000 27.200 ;
        RECT 9.400 27.100 9.800 27.200 ;
        RECT 8.600 26.800 9.800 27.100 ;
        RECT 10.200 26.200 10.500 27.800 ;
        RECT 11.800 27.200 12.100 31.800 ;
        RECT 11.800 26.800 12.200 27.200 ;
        RECT 13.400 26.200 13.700 31.800 ;
        RECT 15.800 29.800 16.200 30.200 ;
        RECT 15.800 29.200 16.100 29.800 ;
        RECT 15.800 28.800 16.200 29.200 ;
        RECT 15.000 28.100 15.400 28.200 ;
        RECT 15.800 28.100 16.200 28.200 ;
        RECT 15.000 27.800 16.200 28.100 ;
        RECT 15.000 26.800 15.400 27.200 ;
        RECT 15.000 26.200 15.300 26.800 ;
        RECT 3.000 25.800 4.100 26.100 ;
        RECT 6.200 25.800 6.600 26.200 ;
        RECT 9.400 25.800 9.800 26.200 ;
        RECT 10.200 25.800 10.600 26.200 ;
        RECT 13.400 25.800 13.800 26.200 ;
        RECT 15.000 25.800 15.400 26.200 ;
        RECT 3.000 24.800 3.400 25.200 ;
        RECT 3.000 24.200 3.300 24.800 ;
        RECT 3.000 23.800 3.400 24.200 ;
        RECT 3.000 14.200 3.300 23.800 ;
        RECT 3.800 15.200 4.100 25.800 ;
        RECT 8.600 24.800 9.000 25.200 ;
        RECT 8.600 24.200 8.900 24.800 ;
        RECT 5.400 24.100 5.800 24.200 ;
        RECT 6.200 24.100 6.600 24.200 ;
        RECT 5.400 23.800 6.600 24.100 ;
        RECT 8.600 23.800 9.000 24.200 ;
        RECT 7.000 22.800 7.400 23.200 ;
        RECT 7.000 22.200 7.300 22.800 ;
        RECT 7.000 21.800 7.400 22.200 ;
        RECT 9.400 19.200 9.700 25.800 ;
        RECT 9.400 18.800 9.800 19.200 ;
        RECT 9.400 17.200 9.700 18.800 ;
        RECT 7.800 16.800 8.200 17.200 ;
        RECT 9.400 16.800 9.800 17.200 ;
        RECT 7.800 16.200 8.100 16.800 ;
        RECT 7.800 15.800 8.200 16.200 ;
        RECT 3.800 14.800 4.200 15.200 ;
        RECT 9.400 14.800 9.800 15.200 ;
        RECT 3.000 13.800 3.400 14.200 ;
        RECT 4.600 14.100 5.000 14.200 ;
        RECT 5.400 14.100 5.800 14.200 ;
        RECT 4.600 13.800 5.800 14.100 ;
        RECT 9.400 13.200 9.700 14.800 ;
        RECT 10.200 13.200 10.500 25.800 ;
        RECT 15.800 25.200 16.100 27.800 ;
        RECT 16.600 27.200 16.900 35.800 ;
        RECT 18.200 34.800 18.600 35.200 ;
        RECT 18.200 34.200 18.500 34.800 ;
        RECT 19.000 34.200 19.300 36.800 ;
        RECT 24.600 35.200 24.900 38.800 ;
        RECT 33.400 38.200 33.700 41.800 ;
        RECT 33.400 37.800 33.800 38.200 ;
        RECT 36.600 37.200 36.900 46.800 ;
        RECT 38.200 45.200 38.500 50.800 ;
        RECT 39.000 47.800 39.400 48.200 ;
        RECT 39.000 46.200 39.300 47.800 ;
        RECT 39.800 47.200 40.100 55.800 ;
        RECT 41.400 55.200 41.700 61.800 ;
        RECT 43.800 57.200 44.100 62.800 ;
        RECT 43.800 56.800 44.200 57.200 ;
        RECT 47.000 56.200 47.300 66.800 ;
        RECT 47.800 66.200 48.100 67.800 ;
        RECT 50.200 66.200 50.500 70.800 ;
        RECT 53.400 68.800 53.800 69.200 ;
        RECT 53.400 68.200 53.700 68.800 ;
        RECT 53.400 67.800 53.800 68.200 ;
        RECT 55.000 67.200 55.300 73.800 ;
        RECT 60.600 72.800 61.000 73.200 ;
        RECT 59.000 72.100 59.400 72.200 ;
        RECT 59.800 72.100 60.200 72.200 ;
        RECT 59.000 71.800 60.200 72.100 ;
        RECT 55.800 70.800 56.200 71.200 ;
        RECT 51.000 66.800 51.400 67.200 ;
        RECT 51.800 66.800 52.200 67.200 ;
        RECT 52.600 67.100 53.000 67.200 ;
        RECT 53.400 67.100 53.800 67.200 ;
        RECT 52.600 66.800 53.800 67.100 ;
        RECT 54.200 66.800 54.600 67.200 ;
        RECT 55.000 66.800 55.400 67.200 ;
        RECT 47.800 65.800 48.200 66.200 ;
        RECT 50.200 65.800 50.600 66.200 ;
        RECT 47.800 65.100 48.200 65.200 ;
        RECT 48.600 65.100 49.000 65.200 ;
        RECT 47.800 64.800 49.000 65.100 ;
        RECT 50.200 64.800 50.600 65.200 ;
        RECT 50.200 64.200 50.500 64.800 ;
        RECT 50.200 63.800 50.600 64.200 ;
        RECT 51.000 60.200 51.300 66.800 ;
        RECT 51.800 61.200 52.100 66.800 ;
        RECT 53.400 61.800 53.800 62.200 ;
        RECT 51.800 60.800 52.200 61.200 ;
        RECT 51.000 59.800 51.400 60.200 ;
        RECT 48.600 58.800 49.000 59.200 ;
        RECT 48.600 58.200 48.900 58.800 ;
        RECT 48.600 57.800 49.000 58.200 ;
        RECT 47.000 55.800 47.400 56.200 ;
        RECT 48.600 56.100 49.000 56.200 ;
        RECT 49.400 56.100 49.800 56.200 ;
        RECT 48.600 55.800 49.800 56.100 ;
        RECT 41.400 54.800 41.800 55.200 ;
        RECT 42.200 54.800 42.600 55.200 ;
        RECT 46.200 55.100 46.600 55.200 ;
        RECT 47.000 55.100 47.400 55.200 ;
        RECT 46.200 54.800 47.400 55.100 ;
        RECT 42.200 54.200 42.500 54.800 ;
        RECT 51.000 54.200 51.300 59.800 ;
        RECT 53.400 56.200 53.700 61.800 ;
        RECT 51.800 56.100 52.200 56.200 ;
        RECT 52.600 56.100 53.000 56.200 ;
        RECT 51.800 55.800 53.000 56.100 ;
        RECT 53.400 55.800 53.800 56.200 ;
        RECT 51.800 55.100 52.200 55.200 ;
        RECT 52.600 55.100 53.000 55.200 ;
        RECT 51.800 54.800 53.000 55.100 ;
        RECT 53.400 54.800 53.800 55.200 ;
        RECT 41.400 53.800 41.800 54.200 ;
        RECT 42.200 53.800 42.600 54.200 ;
        RECT 47.000 53.800 47.400 54.200 ;
        RECT 51.000 53.800 51.400 54.200 ;
        RECT 41.400 51.200 41.700 53.800 ;
        RECT 43.800 52.800 44.200 53.200 ;
        RECT 41.400 50.800 41.800 51.200 ;
        RECT 42.200 48.800 42.600 49.200 ;
        RECT 39.800 46.800 40.200 47.200 ;
        RECT 39.800 46.200 40.100 46.800 ;
        RECT 42.200 46.200 42.500 48.800 ;
        RECT 43.800 47.200 44.100 52.800 ;
        RECT 44.600 51.800 45.000 52.200 ;
        RECT 45.400 51.800 45.800 52.200 ;
        RECT 44.600 50.200 44.900 51.800 ;
        RECT 44.600 49.800 45.000 50.200 ;
        RECT 45.400 47.200 45.700 51.800 ;
        RECT 47.000 49.200 47.300 53.800 ;
        RECT 47.800 52.800 48.200 53.200 ;
        RECT 49.400 53.100 49.800 53.200 ;
        RECT 50.200 53.100 50.600 53.200 ;
        RECT 49.400 52.800 50.600 53.100 ;
        RECT 47.800 49.200 48.100 52.800 ;
        RECT 50.200 51.800 50.600 52.200 ;
        RECT 50.200 49.200 50.500 51.800 ;
        RECT 51.000 50.800 51.400 51.200 ;
        RECT 47.000 48.800 47.400 49.200 ;
        RECT 47.800 48.800 48.200 49.200 ;
        RECT 50.200 48.800 50.600 49.200 ;
        RECT 46.200 47.800 46.600 48.200 ;
        RECT 48.600 47.800 49.000 48.200 ;
        RECT 43.800 46.800 44.200 47.200 ;
        RECT 44.600 46.800 45.000 47.200 ;
        RECT 45.400 46.800 45.800 47.200 ;
        RECT 44.600 46.200 44.900 46.800 ;
        RECT 39.000 45.800 39.400 46.200 ;
        RECT 39.800 45.800 40.200 46.200 ;
        RECT 40.600 45.800 41.000 46.200 ;
        RECT 42.200 45.800 42.600 46.200 ;
        RECT 43.000 45.800 43.400 46.200 ;
        RECT 44.600 45.800 45.000 46.200 ;
        RECT 38.200 44.800 38.600 45.200 ;
        RECT 38.200 42.800 38.600 43.200 ;
        RECT 38.200 39.200 38.500 42.800 ;
        RECT 38.200 38.800 38.600 39.200 ;
        RECT 36.600 36.800 37.000 37.200 ;
        RECT 30.200 36.100 30.600 36.200 ;
        RECT 31.000 36.100 31.400 36.200 ;
        RECT 30.200 35.800 31.400 36.100 ;
        RECT 35.000 35.800 35.400 36.200 ;
        RECT 20.600 35.100 21.000 35.200 ;
        RECT 21.400 35.100 21.800 35.200 ;
        RECT 20.600 34.800 21.800 35.100 ;
        RECT 24.600 34.800 25.000 35.200 ;
        RECT 28.600 35.100 29.000 35.200 ;
        RECT 29.400 35.100 29.800 35.200 ;
        RECT 28.600 34.800 29.800 35.100 ;
        RECT 33.400 35.100 33.800 35.200 ;
        RECT 34.200 35.100 34.600 35.200 ;
        RECT 33.400 34.800 34.600 35.100 ;
        RECT 18.200 33.800 18.600 34.200 ;
        RECT 19.000 33.800 19.400 34.200 ;
        RECT 22.200 33.800 22.600 34.200 ;
        RECT 23.000 34.100 23.400 34.200 ;
        RECT 23.800 34.100 24.200 34.200 ;
        RECT 23.000 33.800 24.200 34.100 ;
        RECT 19.000 33.200 19.300 33.800 ;
        RECT 22.200 33.200 22.500 33.800 ;
        RECT 19.000 32.800 19.400 33.200 ;
        RECT 20.600 32.800 21.000 33.200 ;
        RECT 22.200 32.800 22.600 33.200 ;
        RECT 23.000 33.100 23.400 33.200 ;
        RECT 23.800 33.100 24.200 33.200 ;
        RECT 23.000 32.800 24.200 33.100 ;
        RECT 19.000 32.100 19.400 32.200 ;
        RECT 19.800 32.100 20.200 32.200 ;
        RECT 19.000 31.800 20.200 32.100 ;
        RECT 20.600 31.200 20.900 32.800 ;
        RECT 20.600 30.800 21.000 31.200 ;
        RECT 24.600 28.200 24.900 34.800 ;
        RECT 35.000 34.200 35.300 35.800 ;
        RECT 38.200 34.800 38.600 35.200 ;
        RECT 27.000 33.800 27.400 34.200 ;
        RECT 33.400 33.800 33.800 34.200 ;
        RECT 35.000 34.100 35.400 34.200 ;
        RECT 34.200 33.800 35.400 34.100 ;
        RECT 37.400 33.800 37.800 34.200 ;
        RECT 27.000 32.200 27.300 33.800 ;
        RECT 27.000 31.800 27.400 32.200 ;
        RECT 29.400 31.800 29.800 32.200 ;
        RECT 32.600 31.800 33.000 32.200 ;
        RECT 24.600 27.800 25.000 28.200 ;
        RECT 16.600 26.800 17.000 27.200 ;
        RECT 18.200 27.100 18.600 27.200 ;
        RECT 19.000 27.100 19.400 27.200 ;
        RECT 18.200 26.800 19.400 27.100 ;
        RECT 20.600 27.100 21.000 27.200 ;
        RECT 21.400 27.100 21.800 27.200 ;
        RECT 20.600 26.800 21.800 27.100 ;
        RECT 23.800 27.100 24.200 27.200 ;
        RECT 24.600 27.100 25.000 27.200 ;
        RECT 23.800 26.800 25.000 27.100 ;
        RECT 15.800 24.800 16.200 25.200 ;
        RECT 15.000 23.800 15.400 24.200 ;
        RECT 15.000 17.200 15.300 23.800 ;
        RECT 11.000 16.800 11.400 17.200 ;
        RECT 12.600 16.800 13.000 17.200 ;
        RECT 15.000 16.800 15.400 17.200 ;
        RECT 11.000 16.200 11.300 16.800 ;
        RECT 12.600 16.200 12.900 16.800 ;
        RECT 11.000 15.800 11.400 16.200 ;
        RECT 12.600 15.800 13.000 16.200 ;
        RECT 13.400 15.800 13.800 16.200 ;
        RECT 15.000 15.800 15.400 16.200 ;
        RECT 15.800 15.800 16.200 16.200 ;
        RECT 13.400 15.200 13.700 15.800 ;
        RECT 15.000 15.200 15.300 15.800 ;
        RECT 15.800 15.200 16.100 15.800 ;
        RECT 11.800 15.100 12.200 15.200 ;
        RECT 12.600 15.100 13.000 15.200 ;
        RECT 11.800 14.800 13.000 15.100 ;
        RECT 13.400 14.800 13.800 15.200 ;
        RECT 15.000 14.800 15.400 15.200 ;
        RECT 15.800 14.800 16.200 15.200 ;
        RECT 13.400 13.800 13.800 14.200 ;
        RECT 4.600 13.100 5.000 13.200 ;
        RECT 5.400 13.100 5.800 13.200 ;
        RECT 4.600 12.800 5.800 13.100 ;
        RECT 9.400 12.800 9.800 13.200 ;
        RECT 10.200 12.800 10.600 13.200 ;
        RECT 12.600 12.800 13.000 13.200 ;
        RECT 3.800 10.800 4.200 11.200 ;
        RECT 3.800 9.200 4.100 10.800 ;
        RECT 8.600 9.800 9.000 10.200 ;
        RECT 8.600 9.200 8.900 9.800 ;
        RECT 12.600 9.200 12.900 12.800 ;
        RECT 13.400 10.200 13.700 13.800 ;
        RECT 16.600 12.200 16.900 26.800 ;
        RECT 29.400 26.200 29.700 31.800 ;
        RECT 31.000 28.800 31.400 29.200 ;
        RECT 31.000 28.200 31.300 28.800 ;
        RECT 31.000 27.800 31.400 28.200 ;
        RECT 32.600 27.200 32.900 31.800 ;
        RECT 33.400 29.200 33.700 33.800 ;
        RECT 33.400 28.800 33.800 29.200 ;
        RECT 32.600 26.800 33.000 27.200 ;
        RECT 19.000 26.100 19.400 26.200 ;
        RECT 19.800 26.100 20.200 26.200 ;
        RECT 19.000 25.800 20.200 26.100 ;
        RECT 22.200 26.100 22.600 26.200 ;
        RECT 23.000 26.100 23.400 26.200 ;
        RECT 22.200 25.800 23.400 26.100 ;
        RECT 29.400 25.800 29.800 26.200 ;
        RECT 32.600 26.100 33.000 26.200 ;
        RECT 33.400 26.100 33.800 26.200 ;
        RECT 31.800 25.800 33.800 26.100 ;
        RECT 18.200 25.100 18.600 25.200 ;
        RECT 17.400 24.800 18.600 25.100 ;
        RECT 20.600 25.100 21.000 25.200 ;
        RECT 21.400 25.100 21.800 25.200 ;
        RECT 20.600 24.800 21.800 25.100 ;
        RECT 27.000 25.100 27.400 25.200 ;
        RECT 27.800 25.100 28.200 25.200 ;
        RECT 27.000 24.800 28.200 25.100 ;
        RECT 16.600 11.800 17.000 12.200 ;
        RECT 13.400 9.800 13.800 10.200 ;
        RECT 15.800 9.800 16.200 10.200 ;
        RECT 3.800 8.800 4.200 9.200 ;
        RECT 8.600 8.800 9.000 9.200 ;
        RECT 12.600 8.800 13.000 9.200 ;
        RECT 1.400 7.500 1.800 7.900 ;
        RECT 4.500 7.800 4.900 7.900 ;
        RECT 2.100 7.500 4.900 7.800 ;
        RECT 1.400 7.100 1.700 7.500 ;
        RECT 2.100 7.400 2.500 7.500 ;
        RECT 3.800 7.400 4.200 7.500 ;
        RECT 1.400 6.800 4.200 7.100 ;
        RECT 1.400 5.100 1.700 6.800 ;
        RECT 3.900 6.100 4.200 6.800 ;
        RECT 3.900 5.700 4.300 6.100 ;
        RECT 4.600 5.100 4.900 7.500 ;
        RECT 15.800 7.200 16.100 9.800 ;
        RECT 17.400 9.200 17.700 24.800 ;
        RECT 27.800 24.100 28.200 24.200 ;
        RECT 28.600 24.100 29.000 24.200 ;
        RECT 27.800 23.800 29.000 24.100 ;
        RECT 23.000 23.100 23.400 23.200 ;
        RECT 23.800 23.100 24.200 23.200 ;
        RECT 23.000 22.800 24.200 23.100 ;
        RECT 19.000 16.800 19.400 17.200 ;
        RECT 23.000 16.800 23.400 17.200 ;
        RECT 30.200 16.800 30.600 17.200 ;
        RECT 18.200 15.800 18.600 16.200 ;
        RECT 18.200 15.200 18.500 15.800 ;
        RECT 18.200 14.800 18.600 15.200 ;
        RECT 19.000 14.200 19.300 16.800 ;
        RECT 21.400 15.800 21.800 16.200 ;
        RECT 21.400 15.200 21.700 15.800 ;
        RECT 23.000 15.200 23.300 16.800 ;
        RECT 30.200 16.200 30.500 16.800 ;
        RECT 30.200 15.800 30.600 16.200 ;
        RECT 31.000 15.800 31.400 16.200 ;
        RECT 21.400 14.800 21.800 15.200 ;
        RECT 23.000 14.800 23.400 15.200 ;
        RECT 30.200 14.800 30.600 15.200 ;
        RECT 30.200 14.200 30.500 14.800 ;
        RECT 19.000 13.800 19.400 14.200 ;
        RECT 23.800 13.800 24.200 14.200 ;
        RECT 28.600 13.800 29.000 14.200 ;
        RECT 30.200 13.800 30.600 14.200 ;
        RECT 19.800 12.800 20.200 13.200 ;
        RECT 19.800 12.200 20.100 12.800 ;
        RECT 19.000 11.800 19.400 12.200 ;
        RECT 19.800 11.800 20.200 12.200 ;
        RECT 19.000 9.200 19.300 11.800 ;
        RECT 23.800 11.200 24.100 13.800 ;
        RECT 25.400 12.800 25.800 13.200 ;
        RECT 23.800 10.800 24.200 11.200 ;
        RECT 17.400 8.800 17.800 9.200 ;
        RECT 19.000 8.800 19.400 9.200 ;
        RECT 23.800 8.800 24.200 9.200 ;
        RECT 23.800 7.200 24.100 8.800 ;
        RECT 25.400 7.200 25.700 12.800 ;
        RECT 26.200 11.800 26.600 12.200 ;
        RECT 26.200 10.200 26.500 11.800 ;
        RECT 28.600 11.200 28.900 13.800 ;
        RECT 31.000 11.200 31.300 15.800 ;
        RECT 31.800 15.200 32.100 25.800 ;
        RECT 32.600 24.800 33.000 25.200 ;
        RECT 32.600 24.200 32.900 24.800 ;
        RECT 32.600 23.800 33.000 24.200 ;
        RECT 33.400 23.800 33.800 24.200 ;
        RECT 33.400 23.200 33.700 23.800 ;
        RECT 33.400 22.800 33.800 23.200 ;
        RECT 34.200 21.200 34.500 33.800 ;
        RECT 36.600 32.800 37.000 33.200 ;
        RECT 36.600 32.200 36.900 32.800 ;
        RECT 35.800 31.800 36.200 32.200 ;
        RECT 36.600 31.800 37.000 32.200 ;
        RECT 35.800 28.200 36.100 31.800 ;
        RECT 37.400 31.100 37.700 33.800 ;
        RECT 36.600 30.800 37.700 31.100 ;
        RECT 38.200 31.200 38.500 34.800 ;
        RECT 39.800 32.200 40.100 45.800 ;
        RECT 40.600 45.200 40.900 45.800 ;
        RECT 40.600 44.800 41.000 45.200 ;
        RECT 42.200 35.200 42.500 45.800 ;
        RECT 43.000 45.200 43.300 45.800 ;
        RECT 43.000 44.800 43.400 45.200 ;
        RECT 45.400 40.800 45.800 41.200 ;
        RECT 45.400 39.200 45.700 40.800 ;
        RECT 46.200 39.200 46.500 47.800 ;
        RECT 48.600 47.200 48.900 47.800 ;
        RECT 51.000 47.200 51.300 50.800 ;
        RECT 53.400 50.200 53.700 54.800 ;
        RECT 53.400 49.800 53.800 50.200 ;
        RECT 54.200 49.100 54.500 66.800 ;
        RECT 53.400 48.800 54.500 49.100 ;
        RECT 55.000 66.200 55.300 66.800 ;
        RECT 55.800 66.200 56.100 70.800 ;
        RECT 59.000 67.800 59.400 68.200 ;
        RECT 59.000 67.200 59.300 67.800 ;
        RECT 59.000 66.800 59.400 67.200 ;
        RECT 59.800 66.800 60.200 67.200 ;
        RECT 55.000 65.800 55.400 66.200 ;
        RECT 55.800 65.800 56.200 66.200 ;
        RECT 59.000 65.800 59.400 66.200 ;
        RECT 55.000 56.200 55.300 65.800 ;
        RECT 56.600 65.100 57.000 65.200 ;
        RECT 55.800 64.800 57.000 65.100 ;
        RECT 55.000 55.800 55.400 56.200 ;
        RECT 55.000 49.200 55.300 55.800 ;
        RECT 55.800 49.200 56.100 64.800 ;
        RECT 58.200 61.800 58.600 62.200 ;
        RECT 58.200 55.200 58.500 61.800 ;
        RECT 59.000 59.200 59.300 65.800 ;
        RECT 59.800 63.200 60.100 66.800 ;
        RECT 60.600 66.200 60.900 72.800 ;
        RECT 60.600 65.800 61.000 66.200 ;
        RECT 61.400 64.200 61.700 74.800 ;
        RECT 65.400 74.200 65.700 75.800 ;
        RECT 67.000 74.800 67.400 75.200 ;
        RECT 65.400 73.800 65.800 74.200 ;
        RECT 62.200 72.800 62.600 73.200 ;
        RECT 62.200 72.200 62.500 72.800 ;
        RECT 67.000 72.200 67.300 74.800 ;
        RECT 67.800 73.800 68.200 74.200 ;
        RECT 67.800 73.200 68.100 73.800 ;
        RECT 67.800 72.800 68.200 73.200 ;
        RECT 62.200 71.800 62.600 72.200 ;
        RECT 67.000 71.800 67.400 72.200 ;
        RECT 62.200 68.100 62.600 68.200 ;
        RECT 63.000 68.100 63.400 68.200 ;
        RECT 63.800 68.100 64.200 68.200 ;
        RECT 62.200 67.800 64.200 68.100 ;
        RECT 69.400 67.800 69.800 68.200 ;
        RECT 62.200 66.800 62.600 67.200 ;
        RECT 63.000 66.800 63.400 67.200 ;
        RECT 65.400 67.100 65.800 67.200 ;
        RECT 66.200 67.100 66.600 67.200 ;
        RECT 65.400 66.800 66.600 67.100 ;
        RECT 62.200 66.200 62.500 66.800 ;
        RECT 63.000 66.200 63.300 66.800 ;
        RECT 62.200 65.800 62.600 66.200 ;
        RECT 63.000 65.800 63.400 66.200 ;
        RECT 65.400 66.100 65.800 66.200 ;
        RECT 64.600 65.800 65.800 66.100 ;
        RECT 64.600 65.200 64.900 65.800 ;
        RECT 64.600 64.800 65.000 65.200 ;
        RECT 65.400 64.800 65.800 65.200 ;
        RECT 67.800 65.100 68.200 65.200 ;
        RECT 68.600 65.100 69.000 65.200 ;
        RECT 67.800 64.800 69.000 65.100 ;
        RECT 65.400 64.200 65.700 64.800 ;
        RECT 61.400 63.800 61.800 64.200 ;
        RECT 65.400 63.800 65.800 64.200 ;
        RECT 59.800 62.800 60.200 63.200 ;
        RECT 59.800 61.200 60.100 62.800 ;
        RECT 68.600 61.800 69.000 62.200 ;
        RECT 59.800 60.800 60.200 61.200 ;
        RECT 61.400 60.800 61.800 61.200 ;
        RECT 59.000 58.800 59.400 59.200 ;
        RECT 61.400 55.200 61.700 60.800 ;
        RECT 68.600 59.200 68.900 61.800 ;
        RECT 68.600 58.800 69.000 59.200 ;
        RECT 65.400 56.800 65.800 57.200 ;
        RECT 65.400 56.200 65.700 56.800 ;
        RECT 65.400 55.800 65.800 56.200 ;
        RECT 69.400 55.200 69.700 67.800 ;
        RECT 70.200 66.200 70.500 75.800 ;
        RECT 71.000 75.100 71.400 75.200 ;
        RECT 71.800 75.100 72.200 75.200 ;
        RECT 71.000 74.800 72.200 75.100 ;
        RECT 73.400 75.100 73.800 75.200 ;
        RECT 74.200 75.100 74.600 75.200 ;
        RECT 73.400 74.800 74.600 75.100 ;
        RECT 75.800 75.100 76.200 75.200 ;
        RECT 76.600 75.100 77.000 75.200 ;
        RECT 75.800 74.800 77.000 75.100 ;
        RECT 78.200 74.800 78.600 75.200 ;
        RECT 83.800 74.800 84.200 75.200 ;
        RECT 90.200 75.100 90.600 75.200 ;
        RECT 91.000 75.100 91.400 75.200 ;
        RECT 90.200 74.800 91.400 75.100 ;
        RECT 92.600 74.800 93.000 75.200 ;
        RECT 96.600 74.800 97.000 75.200 ;
        RECT 78.200 74.200 78.500 74.800 ;
        RECT 83.800 74.200 84.100 74.800 ;
        RECT 78.200 73.800 78.600 74.200 ;
        RECT 79.000 73.800 79.400 74.200 ;
        RECT 83.800 73.800 84.200 74.200 ;
        RECT 90.200 73.800 90.600 74.200 ;
        RECT 74.200 72.800 74.600 73.200 ;
        RECT 76.600 72.800 77.000 73.200 ;
        RECT 74.200 72.200 74.500 72.800 ;
        RECT 76.600 72.200 76.900 72.800 ;
        RECT 74.200 71.800 74.600 72.200 ;
        RECT 76.600 71.800 77.000 72.200 ;
        RECT 73.400 69.800 73.800 70.200 ;
        RECT 73.400 69.200 73.700 69.800 ;
        RECT 73.400 68.800 73.800 69.200 ;
        RECT 74.200 67.200 74.500 71.800 ;
        RECT 78.200 71.200 78.500 73.800 ;
        RECT 79.000 73.200 79.300 73.800 ;
        RECT 79.000 72.800 79.400 73.200 ;
        RECT 81.400 72.800 81.800 73.200 ;
        RECT 82.200 72.800 82.600 73.200 ;
        RECT 78.200 70.800 78.600 71.200 ;
        RECT 80.600 70.800 81.000 71.200 ;
        RECT 80.600 68.200 80.900 70.800 ;
        RECT 81.400 69.200 81.700 72.800 ;
        RECT 82.200 72.200 82.500 72.800 ;
        RECT 82.200 71.800 82.600 72.200 ;
        RECT 84.600 70.800 85.000 71.200 ;
        RECT 81.400 68.800 81.800 69.200 ;
        RECT 81.400 68.200 81.700 68.800 ;
        RECT 75.000 67.800 75.400 68.200 ;
        RECT 80.600 67.800 81.000 68.200 ;
        RECT 81.400 67.800 81.800 68.200 ;
        RECT 75.000 67.200 75.300 67.800 ;
        RECT 72.600 66.800 73.000 67.200 ;
        RECT 74.200 66.800 74.600 67.200 ;
        RECT 75.000 66.800 75.400 67.200 ;
        RECT 77.400 67.100 77.800 67.200 ;
        RECT 78.200 67.100 78.600 67.200 ;
        RECT 77.400 66.800 78.600 67.100 ;
        RECT 70.200 65.800 70.600 66.200 ;
        RECT 71.000 65.800 71.400 66.200 ;
        RECT 71.000 65.100 71.300 65.800 ;
        RECT 72.600 65.200 72.900 66.800 ;
        RECT 74.200 66.200 74.500 66.800 ;
        RECT 84.600 66.200 84.900 70.800 ;
        RECT 86.200 69.800 86.600 70.200 ;
        RECT 86.200 68.200 86.500 69.800 ;
        RECT 90.200 69.200 90.500 73.800 ;
        RECT 92.600 69.200 92.900 74.800 ;
        RECT 89.400 68.800 89.800 69.200 ;
        RECT 90.200 68.800 90.600 69.200 ;
        RECT 92.600 68.800 93.000 69.200 ;
        RECT 89.400 68.200 89.700 68.800 ;
        RECT 86.200 67.800 86.600 68.200 ;
        RECT 87.800 67.800 88.200 68.200 ;
        RECT 89.400 67.800 89.800 68.200 ;
        RECT 93.400 67.800 93.800 68.200 ;
        RECT 87.800 67.200 88.100 67.800 ;
        RECT 86.200 67.100 86.600 67.200 ;
        RECT 87.000 67.100 87.400 67.200 ;
        RECT 86.200 66.800 87.400 67.100 ;
        RECT 87.800 66.800 88.200 67.200 ;
        RECT 90.200 67.100 90.600 67.200 ;
        RECT 91.000 67.100 91.400 67.200 ;
        RECT 90.200 66.800 91.400 67.100 ;
        RECT 74.200 65.800 74.600 66.200 ;
        RECT 76.600 65.800 77.000 66.200 ;
        RECT 77.400 65.800 77.800 66.200 ;
        RECT 79.800 65.800 80.200 66.200 ;
        RECT 80.600 65.800 81.000 66.200 ;
        RECT 82.200 65.800 82.600 66.200 ;
        RECT 84.600 65.800 85.000 66.200 ;
        RECT 88.600 66.100 89.000 66.200 ;
        RECT 87.800 65.800 89.000 66.100 ;
        RECT 91.800 65.800 92.200 66.200 ;
        RECT 71.000 64.800 72.100 65.100 ;
        RECT 72.600 64.800 73.000 65.200 ;
        RECT 74.200 65.100 74.600 65.200 ;
        RECT 73.400 64.800 74.600 65.100 ;
        RECT 75.800 64.800 76.200 65.200 ;
        RECT 71.800 64.200 72.100 64.800 ;
        RECT 73.400 64.200 73.700 64.800 ;
        RECT 75.800 64.200 76.100 64.800 ;
        RECT 70.200 63.800 70.600 64.200 ;
        RECT 71.000 63.800 71.400 64.200 ;
        RECT 71.800 63.800 72.200 64.200 ;
        RECT 73.400 63.800 73.800 64.200 ;
        RECT 75.800 63.800 76.200 64.200 ;
        RECT 70.200 63.200 70.500 63.800 ;
        RECT 70.200 62.800 70.600 63.200 ;
        RECT 71.000 61.200 71.300 63.800 ;
        RECT 71.000 60.800 71.400 61.200 ;
        RECT 73.400 59.200 73.700 63.800 ;
        RECT 73.400 58.800 73.800 59.200 ;
        RECT 72.600 56.800 73.000 57.200 ;
        RECT 74.200 57.100 74.600 57.200 ;
        RECT 75.000 57.100 75.400 57.200 ;
        RECT 74.200 56.800 75.400 57.100 ;
        RECT 72.600 56.200 72.900 56.800 ;
        RECT 70.200 55.800 70.600 56.200 ;
        RECT 72.600 55.800 73.000 56.200 ;
        RECT 70.200 55.200 70.500 55.800 ;
        RECT 56.600 55.100 57.000 55.200 ;
        RECT 57.400 55.100 57.800 55.200 ;
        RECT 56.600 54.800 57.800 55.100 ;
        RECT 58.200 54.800 58.600 55.200 ;
        RECT 59.800 54.800 60.200 55.200 ;
        RECT 61.400 54.800 61.800 55.200 ;
        RECT 69.400 54.800 69.800 55.200 ;
        RECT 70.200 54.800 70.600 55.200 ;
        RECT 71.800 54.800 72.200 55.200 ;
        RECT 73.400 54.800 73.800 55.200 ;
        RECT 75.800 54.800 76.200 55.200 ;
        RECT 59.800 54.200 60.100 54.800 ;
        RECT 58.200 54.100 58.600 54.200 ;
        RECT 59.000 54.100 59.400 54.200 ;
        RECT 58.200 53.800 59.400 54.100 ;
        RECT 59.800 53.800 60.200 54.200 ;
        RECT 63.800 53.800 64.200 54.200 ;
        RECT 65.400 53.800 65.800 54.200 ;
        RECT 63.800 53.200 64.100 53.800 ;
        RECT 65.400 53.200 65.700 53.800 ;
        RECT 59.800 53.100 60.200 53.200 ;
        RECT 60.600 53.100 61.000 53.200 ;
        RECT 59.800 52.800 61.000 53.100 ;
        RECT 61.400 53.100 61.800 53.200 ;
        RECT 62.200 53.100 62.600 53.200 ;
        RECT 61.400 52.800 62.600 53.100 ;
        RECT 63.800 52.800 64.200 53.200 ;
        RECT 65.400 52.800 65.800 53.200 ;
        RECT 66.200 52.800 66.600 53.200 ;
        RECT 66.200 52.200 66.500 52.800 ;
        RECT 59.000 51.800 59.400 52.200 ;
        RECT 66.200 51.800 66.600 52.200 ;
        RECT 67.000 51.800 67.400 52.200 ;
        RECT 69.400 52.100 69.700 54.800 ;
        RECT 70.200 54.200 70.500 54.800 ;
        RECT 70.200 53.800 70.600 54.200 ;
        RECT 71.800 53.200 72.100 54.800 ;
        RECT 73.400 54.200 73.700 54.800 ;
        RECT 75.800 54.200 76.100 54.800 ;
        RECT 73.400 53.800 73.800 54.200 ;
        RECT 75.800 53.800 76.200 54.200 ;
        RECT 70.200 53.100 70.600 53.200 ;
        RECT 71.000 53.100 71.400 53.200 ;
        RECT 70.200 52.800 71.400 53.100 ;
        RECT 71.800 52.800 72.200 53.200 ;
        RECT 75.000 52.800 75.400 53.200 ;
        RECT 75.800 53.100 76.200 53.200 ;
        RECT 76.600 53.100 76.900 65.800 ;
        RECT 77.400 65.200 77.700 65.800 ;
        RECT 77.400 64.800 77.800 65.200 ;
        RECT 79.800 60.200 80.100 65.800 ;
        RECT 79.800 59.800 80.200 60.200 ;
        RECT 75.800 52.800 76.900 53.100 ;
        RECT 77.400 58.800 77.800 59.200 ;
        RECT 77.400 55.200 77.700 58.800 ;
        RECT 80.600 56.200 80.900 65.800 ;
        RECT 81.400 60.800 81.800 61.200 ;
        RECT 80.600 55.800 81.000 56.200 ;
        RECT 81.400 55.200 81.700 60.800 ;
        RECT 82.200 59.200 82.500 65.800 ;
        RECT 84.600 64.800 85.000 65.200 ;
        RECT 85.400 64.800 85.800 65.200 ;
        RECT 83.000 64.100 83.400 64.200 ;
        RECT 83.800 64.100 84.200 64.200 ;
        RECT 83.000 63.800 84.200 64.100 ;
        RECT 84.600 63.200 84.900 64.800 ;
        RECT 84.600 62.800 85.000 63.200 ;
        RECT 85.400 62.200 85.700 64.800 ;
        RECT 85.400 61.800 85.800 62.200 ;
        RECT 83.000 59.800 83.400 60.200 ;
        RECT 82.200 58.800 82.600 59.200 ;
        RECT 82.200 55.800 82.600 56.200 ;
        RECT 82.200 55.200 82.500 55.800 ;
        RECT 83.000 55.200 83.300 59.800 ;
        RECT 87.800 59.200 88.100 65.800 ;
        RECT 91.800 65.200 92.100 65.800 ;
        RECT 91.800 64.800 92.200 65.200 ;
        RECT 93.400 62.200 93.700 67.800 ;
        RECT 94.200 66.800 94.600 67.200 ;
        RECT 95.800 66.800 96.200 67.200 ;
        RECT 94.200 65.200 94.500 66.800 ;
        RECT 95.800 65.200 96.100 66.800 ;
        RECT 96.600 66.200 96.900 74.800 ;
        RECT 96.600 65.800 97.000 66.200 ;
        RECT 94.200 64.800 94.600 65.200 ;
        RECT 95.800 64.800 96.200 65.200 ;
        RECT 93.400 61.800 93.800 62.200 ;
        RECT 95.000 61.800 95.400 62.200 ;
        RECT 91.000 59.800 91.400 60.200 ;
        RECT 91.000 59.200 91.300 59.800 ;
        RECT 87.800 58.800 88.200 59.200 ;
        RECT 91.000 58.800 91.400 59.200 ;
        RECT 86.200 56.800 86.600 57.200 ;
        RECT 86.200 56.200 86.500 56.800 ;
        RECT 95.000 56.200 95.300 61.800 ;
        RECT 83.800 56.100 84.200 56.200 ;
        RECT 84.600 56.100 85.000 56.200 ;
        RECT 83.800 55.800 85.000 56.100 ;
        RECT 86.200 55.800 86.600 56.200 ;
        RECT 91.000 55.800 91.400 56.200 ;
        RECT 95.000 55.800 95.400 56.200 ;
        RECT 97.400 55.800 97.800 56.200 ;
        RECT 77.400 54.800 77.800 55.200 ;
        RECT 78.200 55.100 78.600 55.200 ;
        RECT 79.000 55.100 79.400 55.200 ;
        RECT 78.200 54.800 79.400 55.100 ;
        RECT 81.400 54.800 81.800 55.200 ;
        RECT 82.200 54.800 82.600 55.200 ;
        RECT 83.000 54.800 83.400 55.200 ;
        RECT 69.400 51.800 71.300 52.100 ;
        RECT 59.000 50.200 59.300 51.800 ;
        RECT 59.000 49.800 59.400 50.200 ;
        RECT 55.000 48.800 55.400 49.200 ;
        RECT 55.800 48.800 56.200 49.200 ;
        RECT 59.000 48.800 59.400 49.200 ;
        RECT 61.400 48.800 61.800 49.200 ;
        RECT 52.600 47.800 53.000 48.200 ;
        RECT 52.600 47.200 52.900 47.800 ;
        RECT 48.600 46.800 49.000 47.200 ;
        RECT 49.400 47.100 49.800 47.200 ;
        RECT 50.200 47.100 50.600 47.200 ;
        RECT 49.400 46.800 50.600 47.100 ;
        RECT 51.000 46.800 51.400 47.200 ;
        RECT 52.600 46.800 53.000 47.200 ;
        RECT 53.400 46.200 53.700 48.800 ;
        RECT 54.200 48.100 54.600 48.200 ;
        RECT 55.000 48.100 55.400 48.200 ;
        RECT 54.200 47.800 55.400 48.100 ;
        RECT 54.200 46.800 54.600 47.200 ;
        RECT 56.600 46.800 57.000 47.200 ;
        RECT 47.800 46.100 48.200 46.200 ;
        RECT 48.600 46.100 49.000 46.200 ;
        RECT 47.800 45.800 49.000 46.100 ;
        RECT 53.400 45.800 53.800 46.200 ;
        RECT 51.800 45.100 52.200 45.200 ;
        RECT 52.600 45.100 53.000 45.200 ;
        RECT 51.800 44.800 53.000 45.100 ;
        RECT 50.200 41.800 50.600 42.200 ;
        RECT 47.000 39.800 47.400 40.200 ;
        RECT 43.800 39.100 44.200 39.200 ;
        RECT 44.600 39.100 45.000 39.200 ;
        RECT 43.800 38.800 45.000 39.100 ;
        RECT 45.400 38.800 45.800 39.200 ;
        RECT 46.200 38.800 46.600 39.200 ;
        RECT 47.000 37.200 47.300 39.800 ;
        RECT 47.000 36.800 47.400 37.200 ;
        RECT 47.800 36.800 48.200 37.200 ;
        RECT 47.800 35.200 48.100 36.800 ;
        RECT 50.200 36.200 50.500 41.800 ;
        RECT 52.600 37.800 53.000 38.200 ;
        RECT 52.600 37.200 52.900 37.800 ;
        RECT 52.600 36.800 53.000 37.200 ;
        RECT 53.400 36.200 53.700 45.800 ;
        RECT 54.200 44.200 54.500 46.800 ;
        RECT 54.200 43.800 54.600 44.200 ;
        RECT 56.600 42.200 56.900 46.800 ;
        RECT 59.000 46.200 59.300 48.800 ;
        RECT 61.400 47.200 61.700 48.800 ;
        RECT 63.800 47.800 64.200 48.200 ;
        RECT 63.800 47.200 64.100 47.800 ;
        RECT 61.400 46.800 61.800 47.200 ;
        RECT 63.800 46.800 64.200 47.200 ;
        RECT 64.600 46.800 65.000 47.200 ;
        RECT 65.400 46.800 65.800 47.200 ;
        RECT 59.000 45.800 59.400 46.200 ;
        RECT 59.800 46.100 60.200 46.200 ;
        RECT 60.600 46.100 61.000 46.200 ;
        RECT 59.800 45.800 61.000 46.100 ;
        RECT 59.000 44.800 59.400 45.200 ;
        RECT 56.600 41.800 57.000 42.200 ;
        RECT 56.600 38.200 56.900 41.800 ;
        RECT 59.000 40.200 59.300 44.800 ;
        RECT 59.800 44.100 60.200 44.200 ;
        RECT 60.600 44.100 61.000 44.200 ;
        RECT 59.800 43.800 61.000 44.100 ;
        RECT 59.000 39.800 59.400 40.200 ;
        RECT 56.600 37.800 57.000 38.200 ;
        RECT 59.000 37.200 59.300 39.800 ;
        RECT 61.400 39.200 61.700 46.800 ;
        RECT 62.200 46.100 62.600 46.200 ;
        RECT 63.000 46.100 63.400 46.200 ;
        RECT 62.200 45.800 63.400 46.100 ;
        RECT 63.800 45.800 64.200 46.200 ;
        RECT 63.800 45.200 64.100 45.800 ;
        RECT 63.800 44.800 64.200 45.200 ;
        RECT 64.600 44.200 64.900 46.800 ;
        RECT 65.400 46.200 65.700 46.800 ;
        RECT 65.400 45.800 65.800 46.200 ;
        RECT 67.000 45.200 67.300 51.800 ;
        RECT 71.000 49.200 71.300 51.800 ;
        RECT 71.000 48.800 71.400 49.200 ;
        RECT 71.800 47.800 72.200 48.200 ;
        RECT 73.400 47.800 73.800 48.200 ;
        RECT 71.800 47.200 72.100 47.800 ;
        RECT 70.200 46.800 70.600 47.200 ;
        RECT 71.800 46.800 72.200 47.200 ;
        RECT 67.800 46.100 68.200 46.200 ;
        RECT 68.600 46.100 69.000 46.200 ;
        RECT 67.800 45.800 69.000 46.100 ;
        RECT 69.400 45.800 69.800 46.200 ;
        RECT 69.400 45.200 69.700 45.800 ;
        RECT 67.000 44.800 67.400 45.200 ;
        RECT 69.400 44.800 69.800 45.200 ;
        RECT 64.600 43.800 65.000 44.200 ;
        RECT 70.200 41.200 70.500 46.800 ;
        RECT 73.400 46.200 73.700 47.800 ;
        RECT 75.000 47.200 75.300 52.800 ;
        RECT 77.400 48.200 77.700 54.800 ;
        RECT 83.000 54.100 83.400 54.200 ;
        RECT 82.200 53.800 83.400 54.100 ;
        RECT 77.400 47.800 77.800 48.200 ;
        RECT 75.000 47.100 75.400 47.200 ;
        RECT 75.800 47.100 76.200 47.200 ;
        RECT 75.000 46.800 76.200 47.100 ;
        RECT 76.600 47.100 77.000 47.200 ;
        RECT 77.400 47.100 77.800 47.200 ;
        RECT 76.600 46.800 77.800 47.100 ;
        RECT 79.000 46.800 79.400 47.200 ;
        RECT 80.600 47.100 81.000 47.200 ;
        RECT 81.400 47.100 81.800 47.200 ;
        RECT 80.600 46.800 81.800 47.100 ;
        RECT 72.600 45.800 73.000 46.200 ;
        RECT 73.400 45.800 73.800 46.200 ;
        RECT 74.200 45.800 74.600 46.200 ;
        RECT 72.600 45.200 72.900 45.800 ;
        RECT 72.600 44.800 73.000 45.200 ;
        RECT 74.200 44.200 74.500 45.800 ;
        RECT 74.200 43.800 74.600 44.200 ;
        RECT 75.800 44.100 76.200 44.200 ;
        RECT 76.600 44.100 77.000 44.200 ;
        RECT 75.800 43.800 77.000 44.100 ;
        RECT 75.000 42.800 75.400 43.200 ;
        RECT 75.000 42.200 75.300 42.800 ;
        RECT 75.000 41.800 75.400 42.200 ;
        RECT 70.200 40.800 70.600 41.200 ;
        RECT 76.600 40.800 77.000 41.200 ;
        RECT 76.600 39.200 76.900 40.800 ;
        RECT 61.400 38.800 61.800 39.200 ;
        RECT 64.600 39.100 65.000 39.200 ;
        RECT 63.800 38.800 65.000 39.100 ;
        RECT 76.600 38.800 77.000 39.200 ;
        RECT 54.200 36.800 54.600 37.200 ;
        RECT 59.000 36.800 59.400 37.200 ;
        RECT 54.200 36.200 54.500 36.800 ;
        RECT 50.200 35.800 50.600 36.200 ;
        RECT 53.400 35.800 53.800 36.200 ;
        RECT 54.200 35.800 54.600 36.200 ;
        RECT 55.800 35.800 56.200 36.200 ;
        RECT 55.800 35.200 56.100 35.800 ;
        RECT 42.200 34.800 42.600 35.200 ;
        RECT 44.600 34.800 45.000 35.200 ;
        RECT 47.800 34.800 48.200 35.200 ;
        RECT 49.400 35.100 49.800 35.200 ;
        RECT 50.200 35.100 50.600 35.200 ;
        RECT 49.400 34.800 50.600 35.100 ;
        RECT 53.400 35.100 53.800 35.200 ;
        RECT 54.200 35.100 54.600 35.200 ;
        RECT 53.400 34.800 54.600 35.100 ;
        RECT 55.800 34.800 56.200 35.200 ;
        RECT 56.600 35.100 57.000 35.200 ;
        RECT 57.400 35.100 57.800 35.200 ;
        RECT 56.600 34.800 57.800 35.100 ;
        RECT 62.200 34.800 62.600 35.200 ;
        RECT 43.800 33.800 44.200 34.200 ;
        RECT 43.800 33.200 44.100 33.800 ;
        RECT 44.600 33.200 44.900 34.800 ;
        RECT 47.800 33.800 48.200 34.200 ;
        RECT 51.800 34.100 52.200 34.200 ;
        RECT 52.600 34.100 53.000 34.200 ;
        RECT 51.800 33.800 53.000 34.100 ;
        RECT 54.200 34.100 54.600 34.200 ;
        RECT 55.000 34.100 55.400 34.200 ;
        RECT 54.200 33.800 55.400 34.100 ;
        RECT 56.600 33.800 57.000 34.200 ;
        RECT 40.600 33.100 41.000 33.200 ;
        RECT 41.400 33.100 41.800 33.200 ;
        RECT 40.600 32.800 41.800 33.100 ;
        RECT 42.200 33.100 42.600 33.200 ;
        RECT 43.000 33.100 43.400 33.200 ;
        RECT 42.200 32.800 43.400 33.100 ;
        RECT 43.800 32.800 44.200 33.200 ;
        RECT 44.600 32.800 45.000 33.200 ;
        RECT 39.000 31.800 39.400 32.200 ;
        RECT 39.800 31.800 40.200 32.200 ;
        RECT 38.200 30.800 38.600 31.200 ;
        RECT 36.600 30.200 36.900 30.800 ;
        RECT 36.600 29.800 37.000 30.200 ;
        RECT 37.400 29.800 37.800 30.200 ;
        RECT 37.400 29.200 37.700 29.800 ;
        RECT 37.400 28.800 37.800 29.200 ;
        RECT 35.800 27.800 36.200 28.200 ;
        RECT 35.000 26.800 35.400 27.200 ;
        RECT 35.000 26.200 35.300 26.800 ;
        RECT 35.000 25.800 35.400 26.200 ;
        RECT 35.800 25.800 36.200 26.200 ;
        RECT 35.800 25.200 36.100 25.800 ;
        RECT 35.800 24.800 36.200 25.200 ;
        RECT 34.200 20.800 34.600 21.200 ;
        RECT 32.600 19.100 33.000 19.200 ;
        RECT 33.400 19.100 33.800 19.200 ;
        RECT 32.600 18.800 33.800 19.100 ;
        RECT 33.400 16.800 33.800 17.200 ;
        RECT 31.800 14.800 32.200 15.200 ;
        RECT 28.600 10.800 29.000 11.200 ;
        RECT 31.000 10.800 31.400 11.200 ;
        RECT 26.200 9.800 26.600 10.200 ;
        RECT 32.600 9.800 33.000 10.200 ;
        RECT 12.600 6.800 13.000 7.200 ;
        RECT 15.800 6.800 16.200 7.200 ;
        RECT 19.000 6.800 19.400 7.200 ;
        RECT 20.600 6.800 21.000 7.200 ;
        RECT 23.800 6.800 24.200 7.200 ;
        RECT 25.400 6.800 25.800 7.200 ;
        RECT 27.000 7.100 27.400 7.200 ;
        RECT 27.800 7.100 28.200 7.200 ;
        RECT 27.000 6.800 28.200 7.100 ;
        RECT 12.600 6.200 12.900 6.800 ;
        RECT 12.600 5.800 13.000 6.200 ;
        RECT 14.200 6.100 14.600 6.200 ;
        RECT 15.000 6.100 15.400 6.200 ;
        RECT 14.200 5.800 15.400 6.100 ;
        RECT 18.200 5.800 18.600 6.200 ;
        RECT 1.400 4.700 1.800 5.100 ;
        RECT 4.500 4.700 4.900 5.100 ;
        RECT 18.200 5.200 18.500 5.800 ;
        RECT 19.000 5.200 19.300 6.800 ;
        RECT 20.600 5.200 20.900 6.800 ;
        RECT 32.600 6.200 32.900 9.800 ;
        RECT 33.400 7.200 33.700 16.800 ;
        RECT 34.200 15.200 34.500 20.800 ;
        RECT 36.600 19.800 37.000 20.200 ;
        RECT 36.600 16.200 36.900 19.800 ;
        RECT 38.200 17.200 38.500 30.800 ;
        RECT 39.000 28.200 39.300 31.800 ;
        RECT 42.200 30.200 42.500 32.800 ;
        RECT 47.800 32.200 48.100 33.800 ;
        RECT 48.600 32.800 49.000 33.200 ;
        RECT 49.400 32.800 49.800 33.200 ;
        RECT 48.600 32.200 48.900 32.800 ;
        RECT 49.400 32.200 49.700 32.800 ;
        RECT 47.800 31.800 48.200 32.200 ;
        RECT 48.600 31.800 49.000 32.200 ;
        RECT 49.400 31.800 49.800 32.200 ;
        RECT 42.200 29.800 42.600 30.200 ;
        RECT 39.000 27.800 39.400 28.200 ;
        RECT 47.800 27.200 48.100 31.800 ;
        RECT 51.000 30.800 51.400 31.200 ;
        RECT 51.000 28.200 51.300 30.800 ;
        RECT 52.600 30.200 52.900 33.800 ;
        RECT 55.000 31.800 55.400 32.200 ;
        RECT 52.600 29.800 53.000 30.200 ;
        RECT 51.000 27.800 51.400 28.200 ;
        RECT 55.000 27.200 55.300 31.800 ;
        RECT 56.600 30.200 56.900 33.800 ;
        RECT 57.400 30.200 57.700 34.800 ;
        RECT 62.200 34.200 62.500 34.800 ;
        RECT 63.800 34.200 64.100 38.800 ;
        RECT 65.400 35.800 65.800 36.200 ;
        RECT 69.400 36.100 69.800 36.200 ;
        RECT 70.200 36.100 70.600 36.200 ;
        RECT 69.400 35.800 70.600 36.100 ;
        RECT 77.400 36.100 77.700 46.800 ;
        RECT 79.000 46.200 79.300 46.800 ;
        RECT 82.200 46.200 82.500 53.800 ;
        RECT 84.600 53.100 85.000 53.200 ;
        RECT 85.400 53.100 85.800 53.200 ;
        RECT 84.600 52.800 85.800 53.100 ;
        RECT 83.000 48.100 83.400 48.200 ;
        RECT 83.800 48.100 84.200 48.200 ;
        RECT 83.000 47.800 84.200 48.100 ;
        RECT 83.800 46.800 84.200 47.200 ;
        RECT 84.600 47.100 85.000 47.200 ;
        RECT 85.400 47.100 85.800 47.200 ;
        RECT 84.600 46.800 85.800 47.100 ;
        RECT 78.200 45.800 78.600 46.200 ;
        RECT 79.000 45.800 79.400 46.200 ;
        RECT 79.800 45.800 80.200 46.200 ;
        RECT 80.600 45.800 81.000 46.200 ;
        RECT 82.200 46.100 82.600 46.200 ;
        RECT 83.000 46.100 83.400 46.200 ;
        RECT 82.200 45.800 83.400 46.100 ;
        RECT 78.200 40.200 78.500 45.800 ;
        RECT 79.800 45.200 80.100 45.800 ;
        RECT 79.800 44.800 80.200 45.200 ;
        RECT 78.200 39.800 78.600 40.200 ;
        RECT 80.600 37.200 80.900 45.800 ;
        RECT 83.800 44.200 84.100 46.800 ;
        RECT 84.600 46.100 85.000 46.200 ;
        RECT 85.400 46.100 85.800 46.200 ;
        RECT 84.600 45.800 85.800 46.100 ;
        RECT 83.800 43.800 84.200 44.200 ;
        RECT 81.400 39.800 81.800 40.200 ;
        RECT 79.800 36.800 80.200 37.200 ;
        RECT 80.600 36.800 81.000 37.200 ;
        RECT 78.200 36.100 78.600 36.200 ;
        RECT 77.400 35.800 78.600 36.100 ;
        RECT 62.200 33.800 62.600 34.200 ;
        RECT 63.000 33.800 63.400 34.200 ;
        RECT 63.800 33.800 64.200 34.200 ;
        RECT 63.000 33.200 63.300 33.800 ;
        RECT 63.000 32.800 63.400 33.200 ;
        RECT 63.800 33.100 64.200 33.200 ;
        RECT 64.600 33.100 65.000 33.200 ;
        RECT 63.800 32.800 65.000 33.100 ;
        RECT 61.400 31.800 61.800 32.200 ;
        RECT 63.000 31.800 63.400 32.200 ;
        RECT 55.800 29.800 56.200 30.200 ;
        RECT 56.600 29.800 57.000 30.200 ;
        RECT 57.400 29.800 57.800 30.200 ;
        RECT 42.200 27.100 42.600 27.200 ;
        RECT 43.000 27.100 43.400 27.200 ;
        RECT 42.200 26.800 43.400 27.100 ;
        RECT 47.800 26.800 48.200 27.200 ;
        RECT 49.400 26.800 49.800 27.200 ;
        RECT 53.400 26.800 53.800 27.200 ;
        RECT 55.000 26.800 55.400 27.200 ;
        RECT 39.000 25.800 39.400 26.200 ;
        RECT 41.400 26.100 41.800 26.200 ;
        RECT 42.200 26.100 42.600 26.200 ;
        RECT 41.400 25.800 42.600 26.100 ;
        RECT 43.000 25.800 43.400 26.200 ;
        RECT 43.800 25.800 44.200 26.200 ;
        RECT 44.600 26.100 45.000 26.200 ;
        RECT 45.400 26.100 45.800 26.200 ;
        RECT 44.600 25.800 45.800 26.100 ;
        RECT 39.000 24.200 39.300 25.800 ;
        RECT 43.000 25.200 43.300 25.800 ;
        RECT 43.000 24.800 43.400 25.200 ;
        RECT 39.000 23.800 39.400 24.200 ;
        RECT 38.200 16.800 38.600 17.200 ;
        RECT 35.800 16.100 36.200 16.200 ;
        RECT 36.600 16.100 37.000 16.200 ;
        RECT 35.800 15.800 37.000 16.100 ;
        RECT 39.000 15.200 39.300 23.800 ;
        RECT 43.800 22.200 44.100 25.800 ;
        RECT 44.600 24.800 45.000 25.200 ;
        RECT 43.800 21.800 44.200 22.200 ;
        RECT 43.000 18.800 43.400 19.200 ;
        RECT 43.000 15.200 43.300 18.800 ;
        RECT 44.600 15.200 44.900 24.800 ;
        RECT 49.400 24.200 49.700 26.800 ;
        RECT 50.200 25.800 50.600 26.200 ;
        RECT 51.000 26.100 51.400 26.200 ;
        RECT 51.800 26.100 52.200 26.200 ;
        RECT 51.000 25.800 52.200 26.100 ;
        RECT 50.200 25.200 50.500 25.800 ;
        RECT 53.400 25.200 53.700 26.800 ;
        RECT 54.200 25.800 54.600 26.200 ;
        RECT 54.200 25.200 54.500 25.800 ;
        RECT 50.200 24.800 50.600 25.200 ;
        RECT 51.000 24.800 51.400 25.200 ;
        RECT 53.400 24.800 53.800 25.200 ;
        RECT 54.200 24.800 54.600 25.200 ;
        RECT 49.400 23.800 49.800 24.200 ;
        RECT 47.800 22.800 48.200 23.200 ;
        RECT 49.400 23.100 49.800 23.200 ;
        RECT 50.200 23.100 50.600 23.200 ;
        RECT 49.400 22.800 50.600 23.100 ;
        RECT 47.000 16.800 47.400 17.200 ;
        RECT 34.200 14.800 34.600 15.200 ;
        RECT 39.000 14.800 39.400 15.200 ;
        RECT 42.200 14.800 42.600 15.200 ;
        RECT 43.000 14.800 43.400 15.200 ;
        RECT 44.600 14.800 45.000 15.200 ;
        RECT 42.200 14.200 42.500 14.800 ;
        RECT 47.000 14.200 47.300 16.800 ;
        RECT 47.800 15.200 48.100 22.800 ;
        RECT 48.600 16.800 49.000 17.200 ;
        RECT 50.200 16.800 50.600 17.200 ;
        RECT 48.600 16.200 48.900 16.800 ;
        RECT 50.200 16.200 50.500 16.800 ;
        RECT 48.600 15.800 49.000 16.200 ;
        RECT 50.200 15.800 50.600 16.200 ;
        RECT 47.800 14.800 48.200 15.200 ;
        RECT 51.000 15.100 51.300 24.800 ;
        RECT 54.200 20.800 54.600 21.200 ;
        RECT 54.200 15.200 54.500 20.800 ;
        RECT 50.200 14.800 51.300 15.100 ;
        RECT 51.800 15.100 52.200 15.200 ;
        RECT 52.600 15.100 53.000 15.200 ;
        RECT 51.800 14.800 53.000 15.100 ;
        RECT 54.200 14.800 54.600 15.200 ;
        RECT 50.200 14.200 50.500 14.800 ;
        RECT 34.200 13.800 34.600 14.200 ;
        RECT 39.000 13.800 39.400 14.200 ;
        RECT 41.400 13.800 41.800 14.200 ;
        RECT 42.200 13.800 42.600 14.200 ;
        RECT 43.000 13.800 43.400 14.200 ;
        RECT 43.800 13.800 44.200 14.200 ;
        RECT 47.000 13.800 47.400 14.200 ;
        RECT 50.200 13.800 50.600 14.200 ;
        RECT 53.400 13.800 53.800 14.200 ;
        RECT 34.200 10.200 34.500 13.800 ;
        RECT 39.000 13.200 39.300 13.800 ;
        RECT 41.400 13.200 41.700 13.800 ;
        RECT 36.600 12.800 37.000 13.200 ;
        RECT 37.400 12.800 37.800 13.200 ;
        RECT 39.000 12.800 39.400 13.200 ;
        RECT 39.800 12.800 40.200 13.200 ;
        RECT 41.400 12.800 41.800 13.200 ;
        RECT 36.600 12.200 36.900 12.800 ;
        RECT 36.600 11.800 37.000 12.200 ;
        RECT 34.200 9.800 34.600 10.200 ;
        RECT 37.400 9.200 37.700 12.800 ;
        RECT 39.800 12.200 40.100 12.800 ;
        RECT 39.800 11.800 40.200 12.200 ;
        RECT 40.600 12.100 41.000 12.200 ;
        RECT 41.400 12.100 41.800 12.200 ;
        RECT 40.600 11.800 41.800 12.100 ;
        RECT 40.600 10.800 41.000 11.200 ;
        RECT 37.400 8.800 37.800 9.200 ;
        RECT 33.400 6.800 33.800 7.200 ;
        RECT 40.600 6.200 40.900 10.800 ;
        RECT 43.000 9.200 43.300 13.800 ;
        RECT 43.800 12.200 44.100 13.800 ;
        RECT 53.400 13.200 53.700 13.800 ;
        RECT 53.400 12.800 53.800 13.200 ;
        RECT 43.800 11.800 44.200 12.200 ;
        RECT 50.200 9.800 50.600 10.200 ;
        RECT 53.400 9.800 53.800 10.200 ;
        RECT 50.200 9.200 50.500 9.800 ;
        RECT 43.000 8.800 43.400 9.200 ;
        RECT 44.600 9.100 45.000 9.200 ;
        RECT 45.400 9.100 45.800 9.200 ;
        RECT 44.600 8.800 45.800 9.100 ;
        RECT 50.200 8.800 50.600 9.200 ;
        RECT 48.700 7.800 49.100 7.900 ;
        RECT 48.700 7.500 51.500 7.800 ;
        RECT 51.800 7.500 52.200 7.900 ;
        RECT 41.400 6.800 41.800 7.200 ;
        RECT 43.800 7.100 44.200 7.200 ;
        RECT 44.600 7.100 45.000 7.200 ;
        RECT 43.800 6.800 45.000 7.100 ;
        RECT 26.200 6.100 26.600 6.200 ;
        RECT 27.000 6.100 27.400 6.200 ;
        RECT 26.200 5.800 27.400 6.100 ;
        RECT 30.200 6.100 30.600 6.200 ;
        RECT 31.000 6.100 31.400 6.200 ;
        RECT 30.200 5.800 31.400 6.100 ;
        RECT 32.600 5.800 33.000 6.200 ;
        RECT 34.200 5.800 34.600 6.200 ;
        RECT 40.600 5.800 41.000 6.200 ;
        RECT 34.200 5.200 34.500 5.800 ;
        RECT 41.400 5.200 41.700 6.800 ;
        RECT 18.200 4.800 18.600 5.200 ;
        RECT 19.000 4.800 19.400 5.200 ;
        RECT 20.600 4.800 21.000 5.200 ;
        RECT 34.200 4.800 34.600 5.200 ;
        RECT 36.600 5.100 37.000 5.200 ;
        RECT 37.400 5.100 37.800 5.200 ;
        RECT 36.600 4.800 37.800 5.100 ;
        RECT 41.400 4.800 41.800 5.200 ;
        RECT 48.700 5.100 49.000 7.500 ;
        RECT 49.400 7.400 49.800 7.500 ;
        RECT 51.100 7.400 51.500 7.500 ;
        RECT 51.900 7.100 52.200 7.500 ;
        RECT 49.400 6.800 52.200 7.100 ;
        RECT 49.400 6.100 49.700 6.800 ;
        RECT 49.300 5.700 49.700 6.100 ;
        RECT 51.900 5.100 52.200 6.800 ;
        RECT 53.400 6.200 53.700 9.800 ;
        RECT 55.000 8.200 55.300 26.800 ;
        RECT 55.800 26.200 56.100 29.800 ;
        RECT 61.400 29.200 61.700 31.800 ;
        RECT 58.200 29.100 58.600 29.200 ;
        RECT 59.000 29.100 59.400 29.200 ;
        RECT 58.200 28.800 59.400 29.100 ;
        RECT 61.400 28.800 61.800 29.200 ;
        RECT 62.200 28.800 62.600 29.200 ;
        RECT 62.200 28.200 62.500 28.800 ;
        RECT 59.000 28.100 59.400 28.200 ;
        RECT 59.800 28.100 60.200 28.200 ;
        RECT 59.000 27.800 60.200 28.100 ;
        RECT 62.200 27.800 62.600 28.200 ;
        RECT 56.600 26.800 57.000 27.200 ;
        RECT 57.400 26.800 57.800 27.200 ;
        RECT 59.800 27.100 60.200 27.200 ;
        RECT 60.600 27.100 61.000 27.200 ;
        RECT 59.800 26.800 61.000 27.100 ;
        RECT 61.400 27.100 61.800 27.200 ;
        RECT 62.200 27.100 62.600 27.200 ;
        RECT 61.400 26.800 62.600 27.100 ;
        RECT 56.600 26.200 56.900 26.800 ;
        RECT 55.800 25.800 56.200 26.200 ;
        RECT 56.600 25.800 57.000 26.200 ;
        RECT 55.800 16.100 56.200 16.200 ;
        RECT 56.600 16.100 56.900 25.800 ;
        RECT 57.400 19.200 57.700 26.800 ;
        RECT 59.000 26.100 59.400 26.200 ;
        RECT 59.800 26.100 60.200 26.200 ;
        RECT 59.000 25.800 60.200 26.100 ;
        RECT 58.200 21.800 58.600 22.200 ;
        RECT 57.400 18.800 57.800 19.200 ;
        RECT 55.800 15.800 56.900 16.100 ;
        RECT 58.200 14.200 58.500 21.800 ;
        RECT 61.400 18.800 61.800 19.200 ;
        RECT 61.400 18.200 61.700 18.800 ;
        RECT 61.400 17.800 61.800 18.200 ;
        RECT 63.000 16.200 63.300 31.800 ;
        RECT 63.800 26.800 64.200 27.200 ;
        RECT 63.800 26.200 64.100 26.800 ;
        RECT 65.400 26.200 65.700 35.800 ;
        RECT 66.200 34.800 66.600 35.200 ;
        RECT 76.600 34.800 77.000 35.200 ;
        RECT 66.200 34.200 66.500 34.800 ;
        RECT 66.200 33.800 66.600 34.200 ;
        RECT 67.000 33.800 67.400 34.200 ;
        RECT 75.800 33.800 76.200 34.200 ;
        RECT 67.000 33.200 67.300 33.800 ;
        RECT 67.000 32.800 67.400 33.200 ;
        RECT 74.200 31.800 74.600 32.200 ;
        RECT 74.200 30.200 74.500 31.800 ;
        RECT 75.800 31.200 76.100 33.800 ;
        RECT 76.600 33.200 76.900 34.800 ;
        RECT 76.600 32.800 77.000 33.200 ;
        RECT 78.200 33.100 78.600 33.200 ;
        RECT 79.000 33.100 79.400 33.200 ;
        RECT 78.200 32.800 79.400 33.100 ;
        RECT 75.800 30.800 76.200 31.200 ;
        RECT 74.200 29.800 74.600 30.200 ;
        RECT 75.800 29.800 76.200 30.200 ;
        RECT 73.400 29.100 73.800 29.200 ;
        RECT 74.200 29.100 74.600 29.200 ;
        RECT 73.400 28.800 74.600 29.100 ;
        RECT 72.600 27.100 73.000 27.200 ;
        RECT 72.600 26.800 73.700 27.100 ;
        RECT 63.800 25.800 64.200 26.200 ;
        RECT 65.400 25.800 65.800 26.200 ;
        RECT 71.000 26.100 71.400 26.200 ;
        RECT 71.800 26.100 72.200 26.200 ;
        RECT 71.000 25.800 72.200 26.100 ;
        RECT 65.400 25.100 65.800 25.200 ;
        RECT 64.600 24.800 65.800 25.100 ;
        RECT 69.400 25.100 69.800 25.200 ;
        RECT 70.200 25.100 70.600 25.200 ;
        RECT 69.400 24.800 70.600 25.100 ;
        RECT 59.000 15.800 59.400 16.200 ;
        RECT 63.000 15.800 63.400 16.200 ;
        RECT 59.000 15.200 59.300 15.800 ;
        RECT 59.000 14.800 59.400 15.200 ;
        RECT 63.000 14.800 63.400 15.200 ;
        RECT 63.800 14.800 64.200 15.200 ;
        RECT 63.000 14.200 63.300 14.800 ;
        RECT 63.800 14.200 64.100 14.800 ;
        RECT 56.600 14.100 57.000 14.200 ;
        RECT 57.400 14.100 57.800 14.200 ;
        RECT 56.600 13.800 57.800 14.100 ;
        RECT 58.200 13.800 58.600 14.200 ;
        RECT 62.200 14.100 62.600 14.200 ;
        RECT 63.000 14.100 63.400 14.200 ;
        RECT 62.200 13.800 63.400 14.100 ;
        RECT 63.800 13.800 64.200 14.200 ;
        RECT 56.600 12.800 57.000 13.200 ;
        RECT 56.600 12.200 56.900 12.800 ;
        RECT 56.600 11.800 57.000 12.200 ;
        RECT 55.000 7.800 55.400 8.200 ;
        RECT 53.400 5.800 53.800 6.200 ;
        RECT 55.800 6.100 56.200 6.200 ;
        RECT 56.600 6.100 56.900 11.800 ;
        RECT 58.200 10.200 58.500 13.800 ;
        RECT 58.200 9.800 58.600 10.200 ;
        RECT 63.800 9.200 64.100 13.800 ;
        RECT 64.600 9.200 64.900 24.800 ;
        RECT 66.200 21.800 66.600 22.200 ;
        RECT 65.400 19.800 65.800 20.200 ;
        RECT 65.400 16.200 65.700 19.800 ;
        RECT 66.200 16.200 66.500 21.800 ;
        RECT 65.400 15.800 65.800 16.200 ;
        RECT 66.200 15.800 66.600 16.200 ;
        RECT 72.600 15.200 72.900 26.800 ;
        RECT 73.400 25.200 73.700 26.800 ;
        RECT 75.000 26.800 75.400 27.200 ;
        RECT 73.400 24.800 73.800 25.200 ;
        RECT 75.000 24.200 75.300 26.800 ;
        RECT 75.800 25.200 76.100 29.800 ;
        RECT 76.600 27.200 76.900 32.800 ;
        RECT 79.800 29.200 80.100 36.800 ;
        RECT 81.400 35.200 81.700 39.800 ;
        RECT 83.800 36.200 84.100 43.800 ;
        RECT 85.400 41.800 85.800 42.200 ;
        RECT 85.400 39.200 85.700 41.800 ;
        RECT 86.200 41.200 86.500 55.800 ;
        RECT 87.000 55.100 87.400 55.200 ;
        RECT 87.800 55.100 88.200 55.200 ;
        RECT 87.000 54.800 88.200 55.100 ;
        RECT 88.600 53.800 89.000 54.200 ;
        RECT 88.600 53.200 88.900 53.800 ;
        RECT 88.600 52.800 89.000 53.200 ;
        RECT 90.200 50.800 90.600 51.200 ;
        RECT 90.200 49.200 90.500 50.800 ;
        RECT 90.200 48.800 90.600 49.200 ;
        RECT 90.200 47.800 90.600 48.200 ;
        RECT 90.200 46.200 90.500 47.800 ;
        RECT 91.000 47.200 91.300 55.800 ;
        RECT 92.600 54.800 93.000 55.200 ;
        RECT 95.000 55.100 95.400 55.200 ;
        RECT 95.800 55.100 96.200 55.200 ;
        RECT 95.000 54.800 96.200 55.100 ;
        RECT 92.600 51.200 92.900 54.800 ;
        RECT 95.000 53.800 95.400 54.200 ;
        RECT 96.600 53.800 97.000 54.200 ;
        RECT 92.600 50.800 93.000 51.200 ;
        RECT 95.000 48.200 95.300 53.800 ;
        RECT 95.000 47.800 95.400 48.200 ;
        RECT 91.000 46.800 91.400 47.200 ;
        RECT 89.400 45.800 89.800 46.200 ;
        RECT 90.200 45.800 90.600 46.200 ;
        RECT 95.000 45.800 95.400 46.200 ;
        RECT 95.800 45.800 96.200 46.200 ;
        RECT 89.400 45.200 89.700 45.800 ;
        RECT 87.000 44.800 87.400 45.200 ;
        RECT 89.400 44.800 89.800 45.200 ;
        RECT 86.200 40.800 86.600 41.200 ;
        RECT 87.000 39.200 87.300 44.800 ;
        RECT 90.200 43.200 90.500 45.800 ;
        RECT 90.200 42.800 90.600 43.200 ;
        RECT 85.400 38.800 85.800 39.200 ;
        RECT 87.000 38.800 87.400 39.200 ;
        RECT 89.400 37.800 89.800 38.200 ;
        RECT 88.600 36.800 89.000 37.200 ;
        RECT 83.800 35.800 84.200 36.200 ;
        RECT 81.400 34.800 81.800 35.200 ;
        RECT 82.200 34.800 82.600 35.200 ;
        RECT 83.800 34.800 84.200 35.200 ;
        RECT 85.400 35.100 85.800 35.200 ;
        RECT 86.200 35.100 86.600 35.200 ;
        RECT 85.400 34.800 86.600 35.100 ;
        RECT 87.800 34.800 88.200 35.200 ;
        RECT 79.800 28.800 80.200 29.200 ;
        RECT 82.200 28.200 82.500 34.800 ;
        RECT 83.000 33.800 83.400 34.200 ;
        RECT 83.000 33.200 83.300 33.800 ;
        RECT 83.000 32.800 83.400 33.200 ;
        RECT 83.800 28.200 84.100 34.800 ;
        RECT 87.800 34.200 88.100 34.800 ;
        RECT 88.600 34.200 88.900 36.800 ;
        RECT 89.400 35.200 89.700 37.800 ;
        RECT 95.000 37.200 95.300 45.800 ;
        RECT 95.800 38.200 96.100 45.800 ;
        RECT 95.800 37.800 96.200 38.200 ;
        RECT 95.000 36.800 95.400 37.200 ;
        RECT 90.200 35.800 90.600 36.200 ;
        RECT 91.000 36.100 91.400 36.200 ;
        RECT 91.800 36.100 92.200 36.200 ;
        RECT 91.000 35.800 92.200 36.100 ;
        RECT 94.200 36.100 94.600 36.200 ;
        RECT 95.000 36.100 95.400 36.200 ;
        RECT 94.200 35.800 95.400 36.100 ;
        RECT 90.200 35.200 90.500 35.800 ;
        RECT 89.400 34.800 89.800 35.200 ;
        RECT 90.200 34.800 90.600 35.200 ;
        RECT 86.200 33.800 86.600 34.200 ;
        RECT 87.800 33.800 88.200 34.200 ;
        RECT 88.600 33.800 89.000 34.200 ;
        RECT 86.200 32.200 86.500 33.800 ;
        RECT 87.000 32.800 87.400 33.200 ;
        RECT 86.200 31.800 86.600 32.200 ;
        RECT 82.200 27.800 82.600 28.200 ;
        RECT 83.800 27.800 84.200 28.200 ;
        RECT 86.200 27.800 86.600 28.200 ;
        RECT 76.600 26.800 77.000 27.200 ;
        RECT 79.000 26.800 79.400 27.200 ;
        RECT 82.200 27.100 82.600 27.200 ;
        RECT 83.000 27.100 83.400 27.200 ;
        RECT 82.200 26.800 83.400 27.100 ;
        RECT 83.800 26.800 84.200 27.200 ;
        RECT 77.400 25.800 77.800 26.200 ;
        RECT 78.200 25.800 78.600 26.200 ;
        RECT 75.800 24.800 76.200 25.200 ;
        RECT 75.000 23.800 75.400 24.200 ;
        RECT 75.000 22.800 75.400 23.200 ;
        RECT 75.000 19.200 75.300 22.800 ;
        RECT 75.000 18.800 75.400 19.200 ;
        RECT 67.800 14.800 68.200 15.200 ;
        RECT 72.600 14.800 73.000 15.200 ;
        RECT 75.800 14.800 76.200 15.200 ;
        RECT 76.600 14.800 77.000 15.200 ;
        RECT 67.800 13.200 68.100 14.800 ;
        RECT 75.800 14.200 76.100 14.800 ;
        RECT 76.600 14.200 76.900 14.800 ;
        RECT 68.600 13.800 69.000 14.200 ;
        RECT 71.000 14.100 71.400 14.200 ;
        RECT 71.800 14.100 72.200 14.200 ;
        RECT 71.000 13.800 72.200 14.100 ;
        RECT 75.800 13.800 76.200 14.200 ;
        RECT 76.600 13.800 77.000 14.200 ;
        RECT 68.600 13.200 68.900 13.800 ;
        RECT 65.400 12.800 65.800 13.200 ;
        RECT 67.800 12.800 68.200 13.200 ;
        RECT 68.600 12.800 69.000 13.200 ;
        RECT 73.400 13.100 73.800 13.200 ;
        RECT 74.200 13.100 74.600 13.200 ;
        RECT 73.400 12.800 74.600 13.100 ;
        RECT 76.600 12.800 77.000 13.200 ;
        RECT 65.400 12.200 65.700 12.800 ;
        RECT 65.400 11.800 65.800 12.200 ;
        RECT 66.200 12.100 66.600 12.200 ;
        RECT 67.000 12.100 67.400 12.200 ;
        RECT 66.200 11.800 67.400 12.100 ;
        RECT 75.000 11.800 75.400 12.200 ;
        RECT 67.000 10.800 67.400 11.200 ;
        RECT 60.600 9.100 61.000 9.200 ;
        RECT 61.400 9.100 61.800 9.200 ;
        RECT 60.600 8.800 61.800 9.100 ;
        RECT 63.800 8.800 64.200 9.200 ;
        RECT 64.600 8.800 65.000 9.200 ;
        RECT 55.800 5.800 56.900 6.100 ;
        RECT 59.000 7.500 59.400 7.900 ;
        RECT 62.100 7.800 62.500 7.900 ;
        RECT 59.700 7.500 62.500 7.800 ;
        RECT 59.000 7.100 59.300 7.500 ;
        RECT 59.700 7.400 60.100 7.500 ;
        RECT 61.400 7.400 61.800 7.500 ;
        RECT 59.000 6.800 61.800 7.100 ;
        RECT 19.000 4.200 19.300 4.800 ;
        RECT 36.600 4.200 36.900 4.800 ;
        RECT 48.700 4.700 49.100 5.100 ;
        RECT 51.800 4.700 52.200 5.100 ;
        RECT 59.000 5.100 59.300 6.800 ;
        RECT 61.500 6.100 61.800 6.800 ;
        RECT 61.500 5.700 61.900 6.100 ;
        RECT 62.200 5.100 62.500 7.500 ;
        RECT 63.800 7.100 64.200 7.200 ;
        RECT 64.600 7.100 65.000 7.200 ;
        RECT 63.800 6.800 65.000 7.100 ;
        RECT 67.000 6.200 67.300 10.800 ;
        RECT 75.000 9.200 75.300 11.800 ;
        RECT 76.600 9.200 76.900 12.800 ;
        RECT 77.400 12.200 77.700 25.800 ;
        RECT 78.200 14.200 78.500 25.800 ;
        RECT 79.000 24.200 79.300 26.800 ;
        RECT 80.600 25.800 81.000 26.200 ;
        RECT 79.000 23.800 79.400 24.200 ;
        RECT 79.000 16.100 79.400 16.200 ;
        RECT 79.800 16.100 80.200 16.200 ;
        RECT 79.000 15.800 80.200 16.100 ;
        RECT 79.000 15.100 79.400 15.200 ;
        RECT 79.800 15.100 80.200 15.200 ;
        RECT 79.000 14.800 80.200 15.100 ;
        RECT 78.200 13.800 78.600 14.200 ;
        RECT 80.600 13.200 80.900 25.800 ;
        RECT 83.800 16.200 84.100 26.800 ;
        RECT 86.200 26.200 86.500 27.800 ;
        RECT 87.000 27.200 87.300 32.800 ;
        RECT 88.600 27.200 88.900 33.800 ;
        RECT 90.200 32.800 90.600 33.200 ;
        RECT 89.400 27.800 89.800 28.200 ;
        RECT 89.400 27.200 89.700 27.800 ;
        RECT 87.000 26.800 87.400 27.200 ;
        RECT 88.600 26.800 89.000 27.200 ;
        RECT 89.400 26.800 89.800 27.200 ;
        RECT 86.200 25.800 86.600 26.200 ;
        RECT 87.000 24.800 87.400 25.200 ;
        RECT 88.600 25.100 89.000 25.200 ;
        RECT 89.400 25.100 89.800 25.200 ;
        RECT 88.600 24.800 89.800 25.100 ;
        RECT 83.800 15.800 84.200 16.200 ;
        RECT 84.600 16.100 85.000 16.200 ;
        RECT 85.400 16.100 85.800 16.200 ;
        RECT 84.600 15.800 85.800 16.100 ;
        RECT 81.400 15.100 81.800 15.200 ;
        RECT 82.200 15.100 82.600 15.200 ;
        RECT 81.400 14.800 82.600 15.100 ;
        RECT 83.000 14.800 83.400 15.200 ;
        RECT 83.800 14.800 84.200 15.200 ;
        RECT 83.000 14.200 83.300 14.800 ;
        RECT 83.800 14.200 84.100 14.800 ;
        RECT 87.000 14.200 87.300 24.800 ;
        RECT 87.800 23.800 88.200 24.200 ;
        RECT 87.800 23.200 88.100 23.800 ;
        RECT 87.800 22.800 88.200 23.200 ;
        RECT 90.200 19.200 90.500 32.800 ;
        RECT 91.800 31.800 92.200 32.200 ;
        RECT 91.000 27.800 91.400 28.200 ;
        RECT 91.000 27.200 91.300 27.800 ;
        RECT 91.000 26.800 91.400 27.200 ;
        RECT 91.800 26.200 92.100 31.800 ;
        RECT 96.600 28.200 96.900 53.800 ;
        RECT 97.400 49.200 97.700 55.800 ;
        RECT 97.400 48.800 97.800 49.200 ;
        RECT 95.000 27.800 95.400 28.200 ;
        RECT 96.600 27.800 97.000 28.200 ;
        RECT 93.400 26.800 93.800 27.200 ;
        RECT 91.800 25.800 92.200 26.200 ;
        RECT 92.600 21.800 93.000 22.200 ;
        RECT 90.200 18.800 90.600 19.200 ;
        RECT 91.000 17.800 91.400 18.200 ;
        RECT 91.000 17.200 91.300 17.800 ;
        RECT 91.000 16.800 91.400 17.200 ;
        RECT 92.600 16.200 92.900 21.800 ;
        RECT 89.400 15.800 89.800 16.200 ;
        RECT 92.600 15.800 93.000 16.200 ;
        RECT 87.800 15.100 88.200 15.200 ;
        RECT 88.600 15.100 89.000 15.200 ;
        RECT 87.800 14.800 89.000 15.100 ;
        RECT 82.200 13.800 82.600 14.200 ;
        RECT 83.000 13.800 83.400 14.200 ;
        RECT 83.800 13.800 84.200 14.200 ;
        RECT 86.200 13.800 86.600 14.200 ;
        RECT 87.000 14.100 87.400 14.200 ;
        RECT 87.800 14.100 88.200 14.200 ;
        RECT 87.000 13.800 88.200 14.100 ;
        RECT 82.200 13.200 82.500 13.800 ;
        RECT 79.000 12.800 79.400 13.200 ;
        RECT 80.600 12.800 81.000 13.200 ;
        RECT 82.200 12.800 82.600 13.200 ;
        RECT 85.400 12.800 85.800 13.200 ;
        RECT 77.400 11.800 77.800 12.200 ;
        RECT 75.000 8.800 75.400 9.200 ;
        RECT 76.600 8.800 77.000 9.200 ;
        RECT 69.400 7.800 69.800 8.200 ;
        RECT 78.200 7.800 78.600 8.200 ;
        RECT 63.800 6.100 64.200 6.200 ;
        RECT 64.600 6.100 65.000 6.200 ;
        RECT 63.800 5.800 65.000 6.100 ;
        RECT 67.000 5.800 67.400 6.200 ;
        RECT 59.000 4.700 59.400 5.100 ;
        RECT 62.100 4.700 62.500 5.100 ;
        RECT 69.400 5.200 69.700 7.800 ;
        RECT 77.400 6.800 77.800 7.200 ;
        RECT 77.400 6.200 77.700 6.800 ;
        RECT 78.200 6.200 78.500 7.800 ;
        RECT 79.000 7.200 79.300 12.800 ;
        RECT 79.800 12.100 80.200 12.200 ;
        RECT 80.600 12.100 81.000 12.200 ;
        RECT 79.800 11.800 81.000 12.100 ;
        RECT 85.400 9.200 85.700 12.800 ;
        RECT 83.800 9.100 84.200 9.200 ;
        RECT 84.600 9.100 85.000 9.200 ;
        RECT 83.800 8.800 85.000 9.100 ;
        RECT 85.400 8.800 85.800 9.200 ;
        RECT 86.200 8.200 86.500 13.800 ;
        RECT 89.400 13.200 89.700 15.800 ;
        RECT 90.200 15.100 90.600 15.200 ;
        RECT 91.000 15.100 91.400 15.200 ;
        RECT 90.200 14.800 91.400 15.100 ;
        RECT 92.600 14.800 93.000 15.200 ;
        RECT 89.400 12.800 89.800 13.200 ;
        RECT 90.200 8.200 90.500 14.800 ;
        RECT 92.600 14.200 92.900 14.800 ;
        RECT 92.600 13.800 93.000 14.200 ;
        RECT 92.600 12.800 93.000 13.200 ;
        RECT 92.600 12.200 92.900 12.800 ;
        RECT 92.600 11.800 93.000 12.200 ;
        RECT 93.400 9.200 93.700 26.800 ;
        RECT 94.200 25.800 94.600 26.200 ;
        RECT 94.200 25.200 94.500 25.800 ;
        RECT 94.200 24.800 94.600 25.200 ;
        RECT 94.200 15.800 94.600 16.200 ;
        RECT 94.200 14.200 94.500 15.800 ;
        RECT 95.000 15.200 95.300 27.800 ;
        RECT 95.800 27.100 96.200 27.200 ;
        RECT 96.600 27.100 97.000 27.200 ;
        RECT 95.800 26.800 97.000 27.100 ;
        RECT 95.800 26.100 96.200 26.200 ;
        RECT 96.600 26.100 97.000 26.200 ;
        RECT 95.800 25.800 97.000 26.100 ;
        RECT 95.000 14.800 95.400 15.200 ;
        RECT 94.200 13.800 94.600 14.200 ;
        RECT 93.400 8.800 93.800 9.200 ;
        RECT 86.200 7.800 86.600 8.200 ;
        RECT 90.200 7.800 90.600 8.200 ;
        RECT 91.800 7.500 92.200 7.900 ;
        RECT 94.900 7.800 95.300 7.900 ;
        RECT 92.500 7.500 95.300 7.800 ;
        RECT 79.000 6.800 79.400 7.200 ;
        RECT 84.600 6.800 85.000 7.200 ;
        RECT 91.800 7.100 92.100 7.500 ;
        RECT 92.500 7.400 92.900 7.500 ;
        RECT 94.200 7.400 94.600 7.500 ;
        RECT 91.800 6.800 94.600 7.100 ;
        RECT 84.600 6.200 84.900 6.800 ;
        RECT 72.600 5.800 73.000 6.200 ;
        RECT 77.400 5.800 77.800 6.200 ;
        RECT 78.200 6.100 78.600 6.200 ;
        RECT 79.000 6.100 79.400 6.200 ;
        RECT 78.200 5.800 79.400 6.100 ;
        RECT 80.600 5.800 81.000 6.200 ;
        RECT 84.600 5.800 85.000 6.200 ;
        RECT 72.600 5.200 72.900 5.800 ;
        RECT 69.400 4.800 69.800 5.200 ;
        RECT 72.600 4.800 73.000 5.200 ;
        RECT 77.400 4.200 77.700 5.800 ;
        RECT 80.600 5.200 80.900 5.800 ;
        RECT 79.000 5.100 79.400 5.200 ;
        RECT 79.800 5.100 80.200 5.200 ;
        RECT 79.000 4.800 80.200 5.100 ;
        RECT 80.600 4.800 81.000 5.200 ;
        RECT 83.800 4.800 84.200 5.200 ;
        RECT 91.800 5.100 92.100 6.800 ;
        RECT 94.300 6.100 94.600 6.800 ;
        RECT 94.300 5.700 94.700 6.100 ;
        RECT 95.000 5.100 95.300 7.500 ;
        RECT 83.800 4.200 84.100 4.800 ;
        RECT 91.800 4.700 92.200 5.100 ;
        RECT 94.900 4.700 95.300 5.100 ;
        RECT 19.000 3.800 19.400 4.200 ;
        RECT 36.600 3.800 37.000 4.200 ;
        RECT 77.400 3.800 77.800 4.200 ;
        RECT 83.800 3.800 84.200 4.200 ;
      LAYER via2 ;
        RECT 39.000 76.800 39.400 77.200 ;
        RECT 17.400 75.800 17.800 76.200 ;
        RECT 72.600 76.800 73.000 77.200 ;
        RECT 76.600 76.800 77.000 77.200 ;
        RECT 50.200 72.800 50.600 73.200 ;
        RECT 5.400 68.800 5.800 69.200 ;
        RECT 12.600 66.800 13.000 67.200 ;
        RECT 54.200 73.800 54.600 74.200 ;
        RECT 53.400 72.800 53.800 73.200 ;
        RECT 47.800 67.800 48.200 68.200 ;
        RECT 24.600 65.800 25.000 66.200 ;
        RECT 11.000 48.800 11.400 49.200 ;
        RECT 3.800 35.800 4.200 36.200 ;
        RECT 27.800 44.800 28.200 45.200 ;
        RECT 17.400 43.800 17.800 44.200 ;
        RECT 25.400 43.800 25.800 44.200 ;
        RECT 44.600 62.800 45.000 63.200 ;
        RECT 33.400 61.800 33.800 62.200 ;
        RECT 31.800 55.800 32.200 56.200 ;
        RECT 5.400 26.800 5.800 27.200 ;
        RECT 9.400 26.800 9.800 27.200 ;
        RECT 5.400 13.800 5.800 14.200 ;
        RECT 47.000 54.800 47.400 55.200 ;
        RECT 52.600 55.800 53.000 56.200 ;
        RECT 52.600 54.800 53.000 55.200 ;
        RECT 21.400 26.800 21.800 27.200 ;
        RECT 24.600 26.800 25.000 27.200 ;
        RECT 12.600 14.800 13.000 15.200 ;
        RECT 32.600 25.800 33.000 26.200 ;
        RECT 27.800 24.800 28.200 25.200 ;
        RECT 23.800 22.800 24.200 23.200 ;
        RECT 63.000 67.800 63.400 68.200 ;
        RECT 71.800 74.800 72.200 75.200 ;
        RECT 91.000 74.800 91.400 75.200 ;
        RECT 87.000 66.800 87.400 67.200 ;
        RECT 75.000 56.800 75.400 57.200 ;
        RECT 57.400 54.800 57.800 55.200 ;
        RECT 59.000 53.800 59.400 54.200 ;
        RECT 60.600 52.800 61.000 53.200 ;
        RECT 62.200 52.800 62.600 53.200 ;
        RECT 50.200 46.800 50.600 47.200 ;
        RECT 48.600 45.800 49.000 46.200 ;
        RECT 52.600 44.800 53.000 45.200 ;
        RECT 44.600 38.800 45.000 39.200 ;
        RECT 60.600 43.800 61.000 44.200 ;
        RECT 63.000 45.800 63.400 46.200 ;
        RECT 68.600 45.800 69.000 46.200 ;
        RECT 64.600 38.800 65.000 39.200 ;
        RECT 54.200 34.800 54.600 35.200 ;
        RECT 57.400 34.800 57.800 35.200 ;
        RECT 43.000 32.800 43.400 33.200 ;
        RECT 27.800 6.800 28.200 7.200 ;
        RECT 64.600 32.800 65.000 33.200 ;
        RECT 43.000 26.800 43.400 27.200 ;
        RECT 42.200 25.800 42.600 26.200 ;
        RECT 45.400 25.800 45.800 26.200 ;
        RECT 51.800 25.800 52.200 26.200 ;
        RECT 50.200 22.800 50.600 23.200 ;
        RECT 41.400 11.800 41.800 12.200 ;
        RECT 45.400 8.800 45.800 9.200 ;
        RECT 44.600 6.800 45.000 7.200 ;
        RECT 27.000 5.800 27.400 6.200 ;
        RECT 37.400 4.800 37.800 5.200 ;
        RECT 59.000 28.800 59.400 29.200 ;
        RECT 59.800 27.800 60.200 28.200 ;
        RECT 74.200 28.800 74.600 29.200 ;
        RECT 57.400 13.800 57.800 14.200 ;
        RECT 91.800 35.800 92.200 36.200 ;
        RECT 83.000 26.800 83.400 27.200 ;
        RECT 71.800 13.800 72.200 14.200 ;
        RECT 67.000 11.800 67.400 12.200 ;
        RECT 61.400 8.800 61.800 9.200 ;
        RECT 82.200 14.800 82.600 15.200 ;
        RECT 64.600 5.800 65.000 6.200 ;
        RECT 80.600 11.800 81.000 12.200 ;
        RECT 84.600 8.800 85.000 9.200 ;
        RECT 91.000 14.800 91.400 15.200 ;
        RECT 96.600 25.800 97.000 26.200 ;
        RECT 79.000 5.800 79.400 6.200 ;
      LAYER metal3 ;
        RECT 39.800 77.800 40.200 78.200 ;
        RECT 37.400 77.100 37.800 77.200 ;
        RECT 13.400 76.800 37.800 77.100 ;
        RECT 39.000 77.100 39.400 77.200 ;
        RECT 39.800 77.100 40.100 77.800 ;
        RECT 39.000 76.800 40.100 77.100 ;
        RECT 72.600 77.100 73.000 77.200 ;
        RECT 75.800 77.100 76.200 77.200 ;
        RECT 76.600 77.100 77.000 77.200 ;
        RECT 72.600 76.800 77.000 77.100 ;
        RECT 13.400 76.200 13.700 76.800 ;
        RECT 11.800 75.800 12.200 76.200 ;
        RECT 13.400 75.800 13.800 76.200 ;
        RECT 17.400 76.100 17.800 76.200 ;
        RECT 19.000 76.100 19.400 76.200 ;
        RECT 17.400 75.800 19.400 76.100 ;
        RECT 25.400 76.100 25.800 76.200 ;
        RECT 26.200 76.100 26.600 76.200 ;
        RECT 25.400 75.800 26.600 76.100 ;
        RECT 64.600 76.100 65.000 76.200 ;
        RECT 71.000 76.100 71.400 76.200 ;
        RECT 64.600 75.800 71.400 76.100 ;
        RECT 11.800 75.100 12.100 75.800 ;
        RECT 16.600 75.100 17.000 75.200 ;
        RECT 11.800 74.800 17.000 75.100 ;
        RECT 71.800 75.100 72.200 75.200 ;
        RECT 73.400 75.100 73.800 75.200 ;
        RECT 75.800 75.100 76.200 75.200 ;
        RECT 71.800 74.800 76.200 75.100 ;
        RECT 91.000 75.100 91.400 75.200 ;
        RECT 96.600 75.100 97.000 75.200 ;
        RECT 91.000 74.800 97.000 75.100 ;
        RECT 54.200 74.100 54.600 74.200 ;
        RECT 65.400 74.100 65.800 74.200 ;
        RECT 78.200 74.100 78.600 74.200 ;
        RECT 54.200 73.800 78.600 74.100 ;
        RECT 79.000 73.800 79.400 74.200 ;
        RECT 83.800 74.100 84.200 74.200 ;
        RECT 90.200 74.100 90.600 74.200 ;
        RECT 83.800 73.800 90.600 74.100 ;
        RECT 79.000 73.200 79.300 73.800 ;
        RECT 23.800 73.100 24.200 73.200 ;
        RECT 28.600 73.100 29.000 73.200 ;
        RECT 23.800 72.800 29.000 73.100 ;
        RECT 35.800 73.100 36.200 73.200 ;
        RECT 37.400 73.100 37.800 73.200 ;
        RECT 35.800 72.800 37.800 73.100 ;
        RECT 50.200 73.100 50.600 73.200 ;
        RECT 53.400 73.100 53.800 73.200 ;
        RECT 60.600 73.100 61.000 73.200 ;
        RECT 50.200 72.800 61.000 73.100 ;
        RECT 62.200 72.800 62.600 73.200 ;
        RECT 67.800 73.100 68.200 73.200 ;
        RECT 70.200 73.100 70.600 73.200 ;
        RECT 67.800 72.800 70.600 73.100 ;
        RECT 79.000 72.800 79.400 73.200 ;
        RECT 82.200 72.800 82.600 73.200 ;
        RECT 62.200 72.200 62.500 72.800 ;
        RECT 82.200 72.200 82.500 72.800 ;
        RECT 15.800 72.100 16.200 72.200 ;
        RECT 30.200 72.100 30.600 72.200 ;
        RECT 35.800 72.100 36.200 72.200 ;
        RECT 15.800 71.800 36.200 72.100 ;
        RECT 45.400 72.100 45.800 72.200 ;
        RECT 51.000 72.100 51.400 72.200 ;
        RECT 45.400 71.800 51.400 72.100 ;
        RECT 59.000 72.100 59.400 72.200 ;
        RECT 61.400 72.100 61.800 72.200 ;
        RECT 59.000 71.800 61.800 72.100 ;
        RECT 62.200 71.800 62.600 72.200 ;
        RECT 67.000 72.100 67.400 72.200 ;
        RECT 74.200 72.100 74.600 72.200 ;
        RECT 67.000 71.800 74.600 72.100 ;
        RECT 76.600 72.100 77.000 72.200 ;
        RECT 76.600 71.800 81.700 72.100 ;
        RECT 82.200 71.800 82.600 72.200 ;
        RECT 3.800 71.100 4.200 71.200 ;
        RECT 21.400 71.100 21.800 71.200 ;
        RECT 47.000 71.100 47.400 71.200 ;
        RECT 50.200 71.100 50.600 71.200 ;
        RECT 3.800 70.800 50.600 71.100 ;
        RECT 55.800 71.100 56.200 71.200 ;
        RECT 67.000 71.100 67.300 71.800 ;
        RECT 55.800 70.800 67.300 71.100 ;
        RECT 78.200 71.100 78.600 71.200 ;
        RECT 80.600 71.100 81.000 71.200 ;
        RECT 78.200 70.800 81.000 71.100 ;
        RECT 81.400 71.100 81.700 71.800 ;
        RECT 84.600 71.100 85.000 71.200 ;
        RECT 81.400 70.800 85.000 71.100 ;
        RECT 22.200 70.100 22.600 70.200 ;
        RECT 31.000 70.100 31.400 70.200 ;
        RECT 37.400 70.100 37.800 70.200 ;
        RECT 22.200 69.800 37.800 70.100 ;
        RECT 73.400 70.100 73.800 70.200 ;
        RECT 86.200 70.100 86.600 70.200 ;
        RECT 73.400 69.800 86.600 70.100 ;
        RECT 4.600 69.100 5.000 69.200 ;
        RECT 5.400 69.100 5.800 69.200 ;
        RECT 4.600 68.800 5.800 69.100 ;
        RECT 7.000 69.100 7.400 69.200 ;
        RECT 23.800 69.100 24.200 69.200 ;
        RECT 7.000 68.800 24.200 69.100 ;
        RECT 24.600 68.800 25.000 69.200 ;
        RECT 39.000 69.100 39.400 69.200 ;
        RECT 53.400 69.100 53.800 69.200 ;
        RECT 89.400 69.100 89.800 69.200 ;
        RECT 39.000 68.800 53.800 69.100 ;
        RECT 59.000 68.800 89.800 69.100 ;
        RECT 4.600 67.800 5.000 68.200 ;
        RECT 10.200 68.100 10.600 68.200 ;
        RECT 19.000 68.100 19.400 68.200 ;
        RECT 24.600 68.100 24.900 68.800 ;
        RECT 59.000 68.200 59.300 68.800 ;
        RECT 10.200 67.800 24.900 68.100 ;
        RECT 35.000 68.100 35.400 68.200 ;
        RECT 39.000 68.100 39.400 68.200 ;
        RECT 42.200 68.100 42.600 68.200 ;
        RECT 35.000 67.800 42.600 68.100 ;
        RECT 47.800 68.100 48.200 68.200 ;
        RECT 59.000 68.100 59.400 68.200 ;
        RECT 63.000 68.100 63.400 68.200 ;
        RECT 47.800 67.800 59.400 68.100 ;
        RECT 62.200 67.800 63.400 68.100 ;
        RECT 69.400 68.100 69.800 68.200 ;
        RECT 70.200 68.100 70.600 68.200 ;
        RECT 75.000 68.100 75.400 68.200 ;
        RECT 69.400 67.800 75.400 68.100 ;
        RECT 81.400 68.100 81.800 68.200 ;
        RECT 87.800 68.100 88.200 68.200 ;
        RECT 81.400 67.800 88.200 68.100 ;
        RECT 4.600 67.100 4.900 67.800 ;
        RECT 12.600 67.100 13.000 67.200 ;
        RECT 4.600 66.800 13.000 67.100 ;
        RECT 26.200 67.100 26.600 67.200 ;
        RECT 30.200 67.100 30.600 67.200 ;
        RECT 32.600 67.100 33.000 67.200 ;
        RECT 26.200 66.800 33.000 67.100 ;
        RECT 52.600 67.100 53.000 67.200 ;
        RECT 54.200 67.100 54.600 67.200 ;
        RECT 62.200 67.100 62.600 67.200 ;
        RECT 52.600 66.800 62.600 67.100 ;
        RECT 65.400 67.100 65.800 67.200 ;
        RECT 66.200 67.100 66.600 67.200 ;
        RECT 65.400 66.800 66.600 67.100 ;
        RECT 74.200 67.100 74.600 67.200 ;
        RECT 77.400 67.100 77.800 67.200 ;
        RECT 74.200 66.800 77.800 67.100 ;
        RECT 87.000 67.100 87.400 67.200 ;
        RECT 90.200 67.100 90.600 67.200 ;
        RECT 94.200 67.100 94.600 67.200 ;
        RECT 87.000 66.800 94.600 67.100 ;
        RECT 8.600 66.100 9.000 66.200 ;
        RECT 12.600 66.100 13.000 66.200 ;
        RECT 8.600 65.800 13.000 66.100 ;
        RECT 14.200 66.100 14.600 66.200 ;
        RECT 17.400 66.100 17.800 66.200 ;
        RECT 14.200 65.800 17.800 66.100 ;
        RECT 24.600 66.100 25.000 66.200 ;
        RECT 43.800 66.100 44.200 66.200 ;
        RECT 24.600 65.800 44.200 66.100 ;
        RECT 55.000 66.100 55.400 66.200 ;
        RECT 63.000 66.100 63.400 66.200 ;
        RECT 70.200 66.100 70.600 66.200 ;
        RECT 76.600 66.100 77.000 66.200 ;
        RECT 77.400 66.100 77.800 66.200 ;
        RECT 55.000 65.800 77.800 66.100 ;
        RECT 7.000 64.800 7.400 65.200 ;
        RECT 15.000 65.100 15.400 65.200 ;
        RECT 22.200 65.100 22.600 65.200 ;
        RECT 15.000 64.800 22.600 65.100 ;
        RECT 46.200 65.100 46.600 65.200 ;
        RECT 47.800 65.100 48.200 65.200 ;
        RECT 64.600 65.100 65.000 65.200 ;
        RECT 46.200 64.800 48.200 65.100 ;
        RECT 50.200 64.800 65.000 65.100 ;
        RECT 65.400 65.100 65.800 65.200 ;
        RECT 67.800 65.100 68.200 65.200 ;
        RECT 72.600 65.100 73.000 65.200 ;
        RECT 65.400 64.800 73.000 65.100 ;
        RECT 75.800 64.800 76.200 65.200 ;
        RECT 84.600 65.100 85.000 65.200 ;
        RECT 91.800 65.100 92.200 65.200 ;
        RECT 95.800 65.100 96.200 65.200 ;
        RECT 84.600 64.800 96.200 65.100 ;
        RECT 7.000 64.200 7.300 64.800 ;
        RECT 15.000 64.200 15.300 64.800 ;
        RECT 50.200 64.200 50.500 64.800 ;
        RECT 7.000 63.800 7.400 64.200 ;
        RECT 15.000 63.800 15.400 64.200 ;
        RECT 15.800 63.800 16.200 64.200 ;
        RECT 22.200 64.100 22.600 64.200 ;
        RECT 37.400 64.100 37.800 64.200 ;
        RECT 22.200 63.800 37.800 64.100 ;
        RECT 50.200 63.800 50.600 64.200 ;
        RECT 61.400 64.100 61.800 64.200 ;
        RECT 70.200 64.100 70.600 64.200 ;
        RECT 61.400 63.800 70.600 64.100 ;
        RECT 71.800 64.100 72.200 64.200 ;
        RECT 73.400 64.100 73.800 64.200 ;
        RECT 71.800 63.800 73.800 64.100 ;
        RECT 75.800 64.100 76.100 64.800 ;
        RECT 83.000 64.100 83.400 64.200 ;
        RECT 75.800 63.800 83.400 64.100 ;
        RECT 12.600 63.100 13.000 63.200 ;
        RECT 15.800 63.100 16.100 63.800 ;
        RECT 12.600 62.800 16.100 63.100 ;
        RECT 21.400 63.100 21.800 63.200 ;
        RECT 43.000 63.100 43.400 63.200 ;
        RECT 21.400 62.800 43.400 63.100 ;
        RECT 44.600 63.100 45.000 63.200 ;
        RECT 59.800 63.100 60.200 63.200 ;
        RECT 44.600 62.800 60.200 63.100 ;
        RECT 17.400 62.100 17.800 62.200 ;
        RECT 26.200 62.100 26.600 62.200 ;
        RECT 17.400 61.800 26.600 62.100 ;
        RECT 33.400 62.100 33.800 62.200 ;
        RECT 39.800 62.100 40.200 62.200 ;
        RECT 33.400 61.800 40.200 62.100 ;
        RECT 51.000 62.100 51.400 62.200 ;
        RECT 79.000 62.100 79.400 62.200 ;
        RECT 84.600 62.100 85.000 62.200 ;
        RECT 85.400 62.100 85.800 62.200 ;
        RECT 51.000 61.800 85.800 62.100 ;
        RECT 90.200 62.100 90.600 62.200 ;
        RECT 93.400 62.100 93.800 62.200 ;
        RECT 90.200 61.800 93.800 62.100 ;
        RECT 7.800 61.100 8.200 61.200 ;
        RECT 21.400 61.100 21.800 61.200 ;
        RECT 7.800 60.800 21.800 61.100 ;
        RECT 35.000 61.100 35.400 61.200 ;
        RECT 47.800 61.100 48.200 61.200 ;
        RECT 51.800 61.100 52.200 61.200 ;
        RECT 35.000 60.800 52.200 61.100 ;
        RECT 59.800 61.100 60.200 61.200 ;
        RECT 61.400 61.100 61.800 61.200 ;
        RECT 59.800 60.800 61.800 61.100 ;
        RECT 71.000 61.100 71.400 61.200 ;
        RECT 81.400 61.100 81.800 61.200 ;
        RECT 71.000 60.800 81.800 61.100 ;
        RECT 3.800 60.100 4.200 60.200 ;
        RECT 25.400 60.100 25.800 60.200 ;
        RECT 3.800 59.800 25.800 60.100 ;
        RECT 51.000 60.100 51.400 60.200 ;
        RECT 79.800 60.100 80.200 60.200 ;
        RECT 83.000 60.100 83.400 60.200 ;
        RECT 91.000 60.100 91.400 60.200 ;
        RECT 51.000 59.800 91.400 60.100 ;
        RECT 7.000 59.100 7.400 59.200 ;
        RECT 35.000 59.100 35.400 59.200 ;
        RECT 59.000 59.100 59.400 59.200 ;
        RECT 61.400 59.100 61.800 59.200 ;
        RECT 7.000 58.800 35.400 59.100 ;
        RECT 48.600 58.800 61.800 59.100 ;
        RECT 68.600 59.100 69.000 59.200 ;
        RECT 77.400 59.100 77.800 59.200 ;
        RECT 82.200 59.100 82.600 59.200 ;
        RECT 68.600 58.800 82.600 59.100 ;
        RECT 48.600 58.200 48.900 58.800 ;
        RECT 11.800 58.100 12.200 58.200 ;
        RECT 11.800 57.800 34.500 58.100 ;
        RECT 48.600 57.800 49.000 58.200 ;
        RECT 34.200 57.200 34.500 57.800 ;
        RECT 14.200 56.800 14.600 57.200 ;
        RECT 22.200 56.800 22.600 57.200 ;
        RECT 34.200 56.800 34.600 57.200 ;
        RECT 37.400 57.100 37.800 57.200 ;
        RECT 43.800 57.100 44.200 57.200 ;
        RECT 37.400 56.800 44.200 57.100 ;
        RECT 65.400 57.100 65.800 57.200 ;
        RECT 72.600 57.100 73.000 57.200 ;
        RECT 65.400 56.800 73.000 57.100 ;
        RECT 75.000 57.100 75.400 57.200 ;
        RECT 86.200 57.100 86.600 57.200 ;
        RECT 75.000 56.800 86.600 57.100 ;
        RECT 14.200 56.100 14.500 56.800 ;
        RECT 22.200 56.200 22.500 56.800 ;
        RECT 19.800 56.100 20.200 56.200 ;
        RECT 14.200 55.800 20.200 56.100 ;
        RECT 22.200 55.800 22.600 56.200 ;
        RECT 31.800 56.100 32.200 56.200 ;
        RECT 35.000 56.100 35.400 56.200 ;
        RECT 31.800 55.800 35.400 56.100 ;
        RECT 39.800 56.100 40.200 56.200 ;
        RECT 47.000 56.100 47.400 56.200 ;
        RECT 48.600 56.100 49.000 56.200 ;
        RECT 39.800 55.800 49.000 56.100 ;
        RECT 52.600 56.100 53.000 56.200 ;
        RECT 53.400 56.100 53.800 56.200 ;
        RECT 52.600 55.800 53.800 56.100 ;
        RECT 70.200 56.100 70.600 56.200 ;
        RECT 82.200 56.100 82.600 56.200 ;
        RECT 83.800 56.100 84.200 56.200 ;
        RECT 70.200 55.800 84.200 56.100 ;
        RECT 91.000 56.100 91.400 56.200 ;
        RECT 95.000 56.100 95.400 56.200 ;
        RECT 91.000 55.800 95.400 56.100 ;
        RECT 47.000 55.100 47.400 55.200 ;
        RECT 52.600 55.100 53.000 55.200 ;
        RECT 36.600 54.800 42.500 55.100 ;
        RECT 47.000 54.800 53.000 55.100 ;
        RECT 57.400 55.100 57.800 55.200 ;
        RECT 59.800 55.100 60.200 55.200 ;
        RECT 71.800 55.100 72.200 55.200 ;
        RECT 78.200 55.100 78.600 55.200 ;
        RECT 57.400 54.800 78.600 55.100 ;
        RECT 83.000 55.100 83.400 55.200 ;
        RECT 87.000 55.100 87.400 55.200 ;
        RECT 83.000 54.800 87.400 55.100 ;
        RECT 95.000 55.100 95.400 55.200 ;
        RECT 95.800 55.100 96.200 55.200 ;
        RECT 95.000 54.800 96.200 55.100 ;
        RECT 36.600 54.200 36.900 54.800 ;
        RECT 42.200 54.200 42.500 54.800 ;
        RECT 21.400 54.100 21.800 54.200 ;
        RECT 24.600 54.100 25.000 54.200 ;
        RECT 21.400 53.800 25.000 54.100 ;
        RECT 36.600 53.800 37.000 54.200 ;
        RECT 42.200 53.800 42.600 54.200 ;
        RECT 59.000 54.100 59.400 54.200 ;
        RECT 65.400 54.100 65.800 54.200 ;
        RECT 70.200 54.100 70.600 54.200 ;
        RECT 59.000 53.800 70.600 54.100 ;
        RECT 73.400 54.100 73.800 54.200 ;
        RECT 75.800 54.100 76.200 54.200 ;
        RECT 73.400 53.800 76.200 54.100 ;
        RECT 4.600 53.100 5.000 53.200 ;
        RECT 7.000 53.100 7.400 53.200 ;
        RECT 4.600 52.800 7.400 53.100 ;
        RECT 10.200 53.100 10.600 53.200 ;
        RECT 11.000 53.100 11.400 53.200 ;
        RECT 11.800 53.100 12.200 53.200 ;
        RECT 10.200 52.800 12.200 53.100 ;
        RECT 13.400 53.100 13.800 53.200 ;
        RECT 16.600 53.100 17.000 53.200 ;
        RECT 17.400 53.100 17.800 53.200 ;
        RECT 13.400 52.800 17.800 53.100 ;
        RECT 49.400 53.100 49.800 53.200 ;
        RECT 51.800 53.100 52.200 53.200 ;
        RECT 49.400 52.800 52.200 53.100 ;
        RECT 60.600 53.100 61.000 53.200 ;
        RECT 62.200 53.100 62.600 53.200 ;
        RECT 60.600 52.800 62.600 53.100 ;
        RECT 63.800 53.100 64.200 53.200 ;
        RECT 64.600 53.100 65.000 53.200 ;
        RECT 63.800 52.800 65.000 53.100 ;
        RECT 70.200 53.100 70.600 53.200 ;
        RECT 75.000 53.100 75.400 53.200 ;
        RECT 70.200 52.800 75.400 53.100 ;
        RECT 84.600 53.100 85.000 53.200 ;
        RECT 88.600 53.100 89.000 53.200 ;
        RECT 84.600 52.800 89.000 53.100 ;
        RECT 15.800 52.100 16.200 52.200 ;
        RECT 8.600 51.800 16.200 52.100 ;
        RECT 20.600 52.100 21.000 52.200 ;
        RECT 39.000 52.100 39.400 52.200 ;
        RECT 45.400 52.100 45.800 52.200 ;
        RECT 20.600 51.800 45.800 52.100 ;
        RECT 50.200 52.100 50.600 52.200 ;
        RECT 62.200 52.100 62.600 52.200 ;
        RECT 66.200 52.100 66.600 52.200 ;
        RECT 50.200 51.800 66.600 52.100 ;
        RECT 8.600 51.200 8.900 51.800 ;
        RECT 8.600 50.800 9.000 51.200 ;
        RECT 10.200 51.100 10.600 51.200 ;
        RECT 11.000 51.100 11.400 51.200 ;
        RECT 10.200 50.800 11.400 51.100 ;
        RECT 16.600 51.100 17.000 51.200 ;
        RECT 31.000 51.100 31.400 51.200 ;
        RECT 16.600 50.800 31.400 51.100 ;
        RECT 38.200 51.100 38.600 51.200 ;
        RECT 41.400 51.100 41.800 51.200 ;
        RECT 51.000 51.100 51.400 51.200 ;
        RECT 38.200 50.800 51.400 51.100 ;
        RECT 90.200 51.100 90.600 51.200 ;
        RECT 92.600 51.100 93.000 51.200 ;
        RECT 90.200 50.800 93.000 51.100 ;
        RECT 26.200 50.100 26.600 50.200 ;
        RECT 37.400 50.100 37.800 50.200 ;
        RECT 26.200 49.800 37.800 50.100 ;
        RECT 44.600 50.100 45.000 50.200 ;
        RECT 45.400 50.100 45.800 50.200 ;
        RECT 44.600 49.800 45.800 50.100 ;
        RECT 53.400 50.100 53.800 50.200 ;
        RECT 54.200 50.100 54.600 50.200 ;
        RECT 53.400 49.800 54.600 50.100 ;
        RECT 59.000 50.100 59.400 50.200 ;
        RECT 67.000 50.100 67.400 50.200 ;
        RECT 59.000 49.800 67.400 50.100 ;
        RECT 9.400 49.100 9.800 49.200 ;
        RECT 11.000 49.100 11.400 49.200 ;
        RECT 13.400 49.100 13.800 49.200 ;
        RECT 9.400 48.800 13.800 49.100 ;
        RECT 15.800 49.100 16.200 49.200 ;
        RECT 23.800 49.100 24.200 49.200 ;
        RECT 15.800 48.800 24.200 49.100 ;
        RECT 27.000 49.100 27.400 49.200 ;
        RECT 42.200 49.100 42.600 49.200 ;
        RECT 47.800 49.100 48.200 49.200 ;
        RECT 27.000 48.800 48.200 49.100 ;
        RECT 55.000 49.100 55.400 49.200 ;
        RECT 59.000 49.100 59.400 49.200 ;
        RECT 55.000 48.800 59.400 49.100 ;
        RECT 61.400 49.100 61.800 49.200 ;
        RECT 61.400 48.800 88.900 49.100 ;
        RECT 88.600 48.200 88.900 48.800 ;
        RECT 11.000 48.100 11.400 48.200 ;
        RECT 18.200 48.100 18.600 48.200 ;
        RECT 19.800 48.100 20.200 48.200 ;
        RECT 11.000 47.800 20.200 48.100 ;
        RECT 35.800 48.100 36.200 48.200 ;
        RECT 39.000 48.100 39.400 48.200 ;
        RECT 35.800 47.800 39.400 48.100 ;
        RECT 43.800 48.100 44.200 48.200 ;
        RECT 48.600 48.100 49.000 48.200 ;
        RECT 43.800 47.800 49.000 48.100 ;
        RECT 52.600 48.100 53.000 48.200 ;
        RECT 54.200 48.100 54.600 48.200 ;
        RECT 52.600 47.800 54.600 48.100 ;
        RECT 63.800 47.800 64.200 48.200 ;
        RECT 67.000 48.100 67.400 48.200 ;
        RECT 73.400 48.100 73.800 48.200 ;
        RECT 67.000 47.800 73.800 48.100 ;
        RECT 77.400 48.100 77.800 48.200 ;
        RECT 83.000 48.100 83.400 48.200 ;
        RECT 83.800 48.100 84.200 48.200 ;
        RECT 77.400 47.800 84.200 48.100 ;
        RECT 88.600 48.100 89.000 48.200 ;
        RECT 95.000 48.100 95.400 48.200 ;
        RECT 88.600 47.800 95.400 48.100 ;
        RECT 44.600 47.100 45.000 47.200 ;
        RECT 50.200 47.100 50.600 47.200 ;
        RECT 63.000 47.100 63.400 47.200 ;
        RECT 44.600 46.800 63.400 47.100 ;
        RECT 63.800 47.100 64.100 47.800 ;
        RECT 65.400 47.100 65.800 47.200 ;
        RECT 63.800 46.800 65.800 47.100 ;
        RECT 71.800 47.100 72.200 47.200 ;
        RECT 75.000 47.100 75.400 47.200 ;
        RECT 76.600 47.100 77.000 47.200 ;
        RECT 71.800 46.800 77.000 47.100 ;
        RECT 79.000 46.800 79.400 47.200 ;
        RECT 80.600 47.100 81.000 47.200 ;
        RECT 81.400 47.100 81.800 47.200 ;
        RECT 80.600 46.800 81.800 47.100 ;
        RECT 82.200 47.100 82.600 47.200 ;
        RECT 84.600 47.100 85.000 47.200 ;
        RECT 82.200 46.800 85.000 47.100 ;
        RECT 4.600 46.100 5.000 46.200 ;
        RECT 39.800 46.100 40.200 46.200 ;
        RECT 4.600 45.800 40.200 46.100 ;
        RECT 43.000 45.800 43.400 46.200 ;
        RECT 48.600 46.100 49.000 46.200 ;
        RECT 59.800 46.100 60.200 46.200 ;
        RECT 62.200 46.100 62.600 46.200 ;
        RECT 63.000 46.100 63.400 46.200 ;
        RECT 48.600 45.800 60.900 46.100 ;
        RECT 62.200 45.800 63.400 46.100 ;
        RECT 68.600 46.100 69.000 46.200 ;
        RECT 72.600 46.100 73.000 46.200 ;
        RECT 68.600 45.800 73.000 46.100 ;
        RECT 74.200 46.100 74.600 46.200 ;
        RECT 79.000 46.100 79.300 46.800 ;
        RECT 74.200 45.800 79.300 46.100 ;
        RECT 79.800 46.100 80.200 46.200 ;
        RECT 81.400 46.100 81.800 46.200 ;
        RECT 79.800 45.800 81.800 46.100 ;
        RECT 82.200 46.100 82.600 46.200 ;
        RECT 84.600 46.100 85.000 46.200 ;
        RECT 82.200 45.800 85.000 46.100 ;
        RECT 89.400 45.800 89.800 46.200 ;
        RECT 23.800 45.100 24.200 45.200 ;
        RECT 27.800 45.100 28.200 45.200 ;
        RECT 31.800 45.100 32.200 45.200 ;
        RECT 23.800 44.800 32.200 45.100 ;
        RECT 40.600 45.100 41.000 45.200 ;
        RECT 43.000 45.100 43.300 45.800 ;
        RECT 89.400 45.200 89.700 45.800 ;
        RECT 40.600 44.800 43.300 45.100 ;
        RECT 51.800 45.100 52.200 45.200 ;
        RECT 52.600 45.100 53.000 45.200 ;
        RECT 51.800 44.800 53.000 45.100 ;
        RECT 53.400 45.100 53.800 45.200 ;
        RECT 63.800 45.100 64.200 45.200 ;
        RECT 69.400 45.100 69.800 45.200 ;
        RECT 87.000 45.100 87.400 45.200 ;
        RECT 53.400 44.800 87.400 45.100 ;
        RECT 89.400 44.800 89.800 45.200 ;
        RECT 7.000 44.100 7.400 44.200 ;
        RECT 7.800 44.100 8.200 44.200 ;
        RECT 7.000 43.800 8.200 44.100 ;
        RECT 17.400 44.100 17.800 44.200 ;
        RECT 25.400 44.100 25.800 44.200 ;
        RECT 30.200 44.100 30.600 44.200 ;
        RECT 32.600 44.100 33.000 44.200 ;
        RECT 17.400 43.800 33.000 44.100 ;
        RECT 38.200 43.800 38.600 44.200 ;
        RECT 54.200 44.100 54.600 44.200 ;
        RECT 60.600 44.100 61.000 44.200 ;
        RECT 64.600 44.100 65.000 44.200 ;
        RECT 75.800 44.100 76.200 44.200 ;
        RECT 83.800 44.100 84.200 44.200 ;
        RECT 54.200 43.800 84.200 44.100 ;
        RECT 38.200 43.200 38.500 43.800 ;
        RECT 2.200 43.100 2.600 43.200 ;
        RECT 29.400 43.100 29.800 43.200 ;
        RECT 2.200 42.800 29.800 43.100 ;
        RECT 38.200 42.800 38.600 43.200 ;
        RECT 90.200 43.100 90.600 43.200 ;
        RECT 75.000 42.800 90.600 43.100 ;
        RECT 75.000 42.200 75.300 42.800 ;
        RECT 7.000 41.800 7.400 42.200 ;
        RECT 29.400 42.100 29.800 42.200 ;
        RECT 56.600 42.100 57.000 42.200 ;
        RECT 29.400 41.800 57.000 42.100 ;
        RECT 75.000 41.800 75.400 42.200 ;
        RECT 75.800 42.100 76.200 42.200 ;
        RECT 85.400 42.100 85.800 42.200 ;
        RECT 75.800 41.800 85.800 42.100 ;
        RECT 7.000 41.200 7.300 41.800 ;
        RECT 1.400 41.100 1.800 41.200 ;
        RECT 3.800 41.100 4.200 41.200 ;
        RECT 1.400 40.800 4.200 41.100 ;
        RECT 7.000 40.800 7.400 41.200 ;
        RECT 45.400 41.100 45.800 41.200 ;
        RECT 70.200 41.100 70.600 41.200 ;
        RECT 45.400 40.800 70.600 41.100 ;
        RECT 76.600 41.100 77.000 41.200 ;
        RECT 86.200 41.100 86.600 41.200 ;
        RECT 76.600 40.800 86.600 41.100 ;
        RECT 47.000 40.100 47.400 40.200 ;
        RECT 59.000 40.100 59.400 40.200 ;
        RECT 47.000 39.800 59.400 40.100 ;
        RECT 78.200 40.100 78.600 40.200 ;
        RECT 81.400 40.100 81.800 40.200 ;
        RECT 78.200 39.800 81.800 40.100 ;
        RECT 8.600 39.100 9.000 39.200 ;
        RECT 24.600 39.100 25.000 39.200 ;
        RECT 8.600 38.800 25.000 39.100 ;
        RECT 44.600 39.100 45.000 39.200 ;
        RECT 46.200 39.100 46.600 39.200 ;
        RECT 61.400 39.100 61.800 39.200 ;
        RECT 44.600 38.800 61.800 39.100 ;
        RECT 63.800 39.100 64.200 39.200 ;
        RECT 64.600 39.100 65.000 39.200 ;
        RECT 63.800 38.800 65.000 39.100 ;
        RECT 20.600 38.100 21.000 38.200 ;
        RECT 23.000 38.100 23.400 38.200 ;
        RECT 20.600 37.800 23.400 38.100 ;
        RECT 23.800 38.100 24.200 38.200 ;
        RECT 33.400 38.100 33.800 38.200 ;
        RECT 23.800 37.800 33.800 38.100 ;
        RECT 52.600 37.800 53.000 38.200 ;
        RECT 53.400 38.100 53.800 38.200 ;
        RECT 56.600 38.100 57.000 38.200 ;
        RECT 53.400 37.800 57.000 38.100 ;
        RECT 89.400 38.100 89.800 38.200 ;
        RECT 95.000 38.100 95.400 38.200 ;
        RECT 95.800 38.100 96.200 38.200 ;
        RECT 89.400 37.800 96.200 38.100 ;
        RECT 10.200 37.100 10.600 37.200 ;
        RECT 11.800 37.100 12.200 37.200 ;
        RECT 19.000 37.100 19.400 37.200 ;
        RECT 36.600 37.100 37.000 37.200 ;
        RECT 10.200 36.800 37.000 37.100 ;
        RECT 47.000 37.100 47.400 37.200 ;
        RECT 47.800 37.100 48.200 37.200 ;
        RECT 47.000 36.800 48.200 37.100 ;
        RECT 52.600 37.100 52.900 37.800 ;
        RECT 54.200 37.100 54.600 37.200 ;
        RECT 52.600 36.800 54.600 37.100 ;
        RECT 59.000 37.100 59.400 37.200 ;
        RECT 79.800 37.100 80.200 37.200 ;
        RECT 59.000 36.800 80.200 37.100 ;
        RECT 88.600 37.100 89.000 37.200 ;
        RECT 95.000 37.100 95.400 37.200 ;
        RECT 88.600 36.800 95.400 37.100 ;
        RECT 3.800 36.100 4.200 36.200 ;
        RECT 5.400 36.100 5.800 36.200 ;
        RECT 3.800 35.800 5.800 36.100 ;
        RECT 9.400 36.100 9.800 36.200 ;
        RECT 14.200 36.100 14.600 36.200 ;
        RECT 9.400 35.800 14.600 36.100 ;
        RECT 16.600 36.100 17.000 36.200 ;
        RECT 30.200 36.100 30.600 36.200 ;
        RECT 35.000 36.100 35.400 36.200 ;
        RECT 16.600 35.800 35.400 36.100 ;
        RECT 43.000 36.100 43.400 36.200 ;
        RECT 50.200 36.100 50.600 36.200 ;
        RECT 43.000 35.800 50.600 36.100 ;
        RECT 53.400 36.100 53.800 36.200 ;
        RECT 55.800 36.100 56.200 36.200 ;
        RECT 65.400 36.100 65.800 36.200 ;
        RECT 53.400 35.800 65.800 36.100 ;
        RECT 67.000 36.100 67.400 36.200 ;
        RECT 69.400 36.100 69.800 36.200 ;
        RECT 67.000 35.800 69.800 36.100 ;
        RECT 90.200 35.800 90.600 36.200 ;
        RECT 91.800 36.100 92.200 36.200 ;
        RECT 94.200 36.100 94.600 36.200 ;
        RECT 91.800 35.800 94.600 36.100 ;
        RECT 3.800 35.100 4.200 35.200 ;
        RECT 7.800 35.100 8.200 35.200 ;
        RECT 3.800 34.800 8.200 35.100 ;
        RECT 13.400 35.100 13.800 35.200 ;
        RECT 14.200 35.100 14.600 35.200 ;
        RECT 13.400 34.800 14.600 35.100 ;
        RECT 18.200 35.100 18.600 35.200 ;
        RECT 20.600 35.100 21.000 35.200 ;
        RECT 18.200 34.800 21.000 35.100 ;
        RECT 28.600 35.100 29.000 35.200 ;
        RECT 33.400 35.100 33.800 35.200 ;
        RECT 28.600 34.800 33.800 35.100 ;
        RECT 42.200 35.100 42.600 35.200 ;
        RECT 49.400 35.100 49.800 35.200 ;
        RECT 50.200 35.100 50.600 35.200 ;
        RECT 42.200 34.800 50.600 35.100 ;
        RECT 54.200 35.100 54.600 35.200 ;
        RECT 57.400 35.100 57.800 35.200 ;
        RECT 54.200 34.800 57.800 35.100 ;
        RECT 83.000 35.100 83.400 35.200 ;
        RECT 83.800 35.100 84.200 35.200 ;
        RECT 83.000 34.800 84.200 35.100 ;
        RECT 85.400 35.100 85.800 35.200 ;
        RECT 87.800 35.100 88.200 35.200 ;
        RECT 90.200 35.100 90.500 35.800 ;
        RECT 85.400 34.800 90.500 35.100 ;
        RECT 23.000 34.100 23.400 34.200 ;
        RECT 43.800 34.100 44.200 34.200 ;
        RECT 23.000 33.800 44.200 34.100 ;
        RECT 47.800 34.100 48.200 34.200 ;
        RECT 51.800 34.100 52.200 34.200 ;
        RECT 47.800 33.800 52.200 34.100 ;
        RECT 54.200 34.100 54.600 34.200 ;
        RECT 62.200 34.100 62.600 34.200 ;
        RECT 54.200 33.800 62.600 34.100 ;
        RECT 66.200 34.100 66.600 34.200 ;
        RECT 70.200 34.100 70.600 34.200 ;
        RECT 66.200 33.800 70.600 34.100 ;
        RECT 0.600 33.100 1.000 33.200 ;
        RECT 9.400 33.100 9.800 33.200 ;
        RECT 0.600 32.800 9.800 33.100 ;
        RECT 19.000 33.100 19.400 33.200 ;
        RECT 22.200 33.100 22.600 33.200 ;
        RECT 19.000 32.800 22.600 33.100 ;
        RECT 23.000 33.100 23.400 33.200 ;
        RECT 24.600 33.100 25.000 33.200 ;
        RECT 23.000 32.800 25.000 33.100 ;
        RECT 40.600 33.100 41.000 33.200 ;
        RECT 41.400 33.100 41.800 33.200 ;
        RECT 40.600 32.800 41.800 33.100 ;
        RECT 43.000 33.100 43.400 33.200 ;
        RECT 44.600 33.100 45.000 33.200 ;
        RECT 63.000 33.100 63.400 33.200 ;
        RECT 43.000 32.800 45.000 33.100 ;
        RECT 48.600 32.800 63.400 33.100 ;
        RECT 64.600 33.100 65.000 33.200 ;
        RECT 67.000 33.100 67.400 33.200 ;
        RECT 64.600 32.800 67.400 33.100 ;
        RECT 76.600 33.100 77.000 33.200 ;
        RECT 78.200 33.100 78.600 33.200 ;
        RECT 76.600 32.800 78.600 33.100 ;
        RECT 82.200 33.100 82.600 33.200 ;
        RECT 83.000 33.100 83.400 33.200 ;
        RECT 87.000 33.100 87.400 33.200 ;
        RECT 82.200 32.800 87.400 33.100 ;
        RECT 89.400 33.100 89.800 33.200 ;
        RECT 90.200 33.100 90.600 33.200 ;
        RECT 89.400 32.800 90.600 33.100 ;
        RECT 48.600 32.200 48.900 32.800 ;
        RECT 19.000 32.100 19.400 32.200 ;
        RECT 27.000 32.100 27.400 32.200 ;
        RECT 29.400 32.100 29.800 32.200 ;
        RECT 19.000 31.800 29.800 32.100 ;
        RECT 36.600 32.100 37.000 32.200 ;
        RECT 39.000 32.100 39.400 32.200 ;
        RECT 36.600 31.800 39.400 32.100 ;
        RECT 39.800 32.100 40.200 32.200 ;
        RECT 47.800 32.100 48.200 32.200 ;
        RECT 39.800 31.800 48.200 32.100 ;
        RECT 48.600 31.800 49.000 32.200 ;
        RECT 49.400 32.100 49.800 32.200 ;
        RECT 55.000 32.100 55.400 32.200 ;
        RECT 49.400 31.800 55.400 32.100 ;
        RECT 61.400 32.100 61.800 32.200 ;
        RECT 86.200 32.100 86.600 32.200 ;
        RECT 91.800 32.100 92.200 32.200 ;
        RECT 61.400 31.800 92.200 32.100 ;
        RECT 6.200 31.100 6.600 31.200 ;
        RECT 19.000 31.100 19.400 31.200 ;
        RECT 20.600 31.100 21.000 31.200 ;
        RECT 6.200 30.800 21.000 31.100 ;
        RECT 38.200 31.100 38.600 31.200 ;
        RECT 51.000 31.100 51.400 31.200 ;
        RECT 38.200 30.800 51.400 31.100 ;
        RECT 72.600 31.100 73.000 31.200 ;
        RECT 75.800 31.100 76.200 31.200 ;
        RECT 72.600 30.800 76.200 31.100 ;
        RECT 4.600 30.100 5.000 30.200 ;
        RECT 6.200 30.100 6.600 30.200 ;
        RECT 4.600 29.800 6.600 30.100 ;
        RECT 15.800 30.100 16.200 30.200 ;
        RECT 36.600 30.100 37.000 30.200 ;
        RECT 15.800 29.800 37.000 30.100 ;
        RECT 37.400 30.100 37.800 30.200 ;
        RECT 42.200 30.100 42.600 30.200 ;
        RECT 37.400 29.800 42.600 30.100 ;
        RECT 52.600 30.100 53.000 30.200 ;
        RECT 55.800 30.100 56.200 30.200 ;
        RECT 52.600 29.800 56.200 30.100 ;
        RECT 56.600 29.800 57.000 30.200 ;
        RECT 57.400 30.100 57.800 30.200 ;
        RECT 62.200 30.100 62.600 30.200 ;
        RECT 57.400 29.800 62.600 30.100 ;
        RECT 70.200 30.100 70.600 30.200 ;
        RECT 74.200 30.100 74.600 30.200 ;
        RECT 75.800 30.100 76.200 30.200 ;
        RECT 70.200 29.800 76.200 30.100 ;
        RECT 56.600 29.200 56.900 29.800 ;
        RECT 31.000 29.100 31.400 29.200 ;
        RECT 43.000 29.100 43.400 29.200 ;
        RECT 31.000 28.800 43.400 29.100 ;
        RECT 56.600 28.800 57.000 29.200 ;
        RECT 59.000 29.100 59.400 29.200 ;
        RECT 59.800 29.100 60.200 29.200 ;
        RECT 58.200 28.800 60.200 29.100 ;
        RECT 62.200 29.100 62.600 29.200 ;
        RECT 63.000 29.100 63.400 29.200 ;
        RECT 74.200 29.100 74.600 29.200 ;
        RECT 62.200 28.800 74.600 29.100 ;
        RECT 10.200 28.100 10.600 28.200 ;
        RECT 15.000 28.100 15.400 28.200 ;
        RECT 10.200 27.800 15.400 28.100 ;
        RECT 35.800 28.100 36.200 28.200 ;
        RECT 42.200 28.100 42.600 28.200 ;
        RECT 35.800 27.800 42.600 28.100 ;
        RECT 43.000 27.800 43.400 28.200 ;
        RECT 44.600 28.100 45.000 28.200 ;
        RECT 59.800 28.100 60.200 28.200 ;
        RECT 82.200 28.100 82.600 28.200 ;
        RECT 86.200 28.100 86.600 28.200 ;
        RECT 89.400 28.100 89.800 28.200 ;
        RECT 44.600 27.800 89.800 28.100 ;
        RECT 91.000 27.800 91.400 28.200 ;
        RECT 95.000 28.100 95.400 28.200 ;
        RECT 96.600 28.100 97.000 28.200 ;
        RECT 95.000 27.800 97.000 28.100 ;
        RECT 43.000 27.200 43.300 27.800 ;
        RECT 5.400 27.100 5.800 27.200 ;
        RECT 9.400 27.100 9.800 27.200 ;
        RECT 5.400 26.800 9.800 27.100 ;
        RECT 14.200 27.100 14.600 27.200 ;
        RECT 15.000 27.100 15.400 27.200 ;
        RECT 14.200 26.800 15.400 27.100 ;
        RECT 18.200 27.100 18.600 27.200 ;
        RECT 19.800 27.100 20.200 27.200 ;
        RECT 18.200 26.800 20.200 27.100 ;
        RECT 21.400 27.100 21.800 27.200 ;
        RECT 23.800 27.100 24.200 27.200 ;
        RECT 24.600 27.100 25.000 27.200 ;
        RECT 21.400 26.800 25.000 27.100 ;
        RECT 32.600 27.100 33.000 27.200 ;
        RECT 38.200 27.100 38.600 27.200 ;
        RECT 32.600 26.800 38.600 27.100 ;
        RECT 43.000 26.800 43.400 27.200 ;
        RECT 56.600 26.800 57.000 27.200 ;
        RECT 59.800 27.100 60.200 27.200 ;
        RECT 60.600 27.100 61.000 27.200 ;
        RECT 59.800 26.800 61.000 27.100 ;
        RECT 61.400 27.100 61.800 27.200 ;
        RECT 62.200 27.100 62.600 27.200 ;
        RECT 61.400 26.800 62.600 27.100 ;
        RECT 63.800 26.800 64.200 27.200 ;
        RECT 83.000 27.100 83.400 27.200 ;
        RECT 88.600 27.100 89.000 27.200 ;
        RECT 91.000 27.100 91.300 27.800 ;
        RECT 93.400 27.100 93.800 27.200 ;
        RECT 95.800 27.100 96.200 27.200 ;
        RECT 83.000 26.800 96.200 27.100 ;
        RECT 7.800 26.100 8.200 26.200 ;
        RECT 9.400 26.100 9.800 26.200 ;
        RECT 7.800 25.800 9.800 26.100 ;
        RECT 13.400 26.100 13.800 26.200 ;
        RECT 19.000 26.100 19.400 26.200 ;
        RECT 22.200 26.100 22.600 26.200 ;
        RECT 13.400 25.800 22.600 26.100 ;
        RECT 32.600 26.100 33.000 26.200 ;
        RECT 35.000 26.100 35.400 26.200 ;
        RECT 39.000 26.100 39.400 26.200 ;
        RECT 32.600 25.800 39.400 26.100 ;
        RECT 42.200 26.100 42.600 26.200 ;
        RECT 45.400 26.100 45.800 26.200 ;
        RECT 42.200 25.800 45.800 26.100 ;
        RECT 47.800 26.100 48.200 26.200 ;
        RECT 51.800 26.100 52.200 26.200 ;
        RECT 56.600 26.100 56.900 26.800 ;
        RECT 47.800 25.800 50.500 26.100 ;
        RECT 51.800 25.800 56.900 26.100 ;
        RECT 59.000 26.100 59.400 26.200 ;
        RECT 59.800 26.100 60.200 26.200 ;
        RECT 59.000 25.800 60.200 26.100 ;
        RECT 61.400 26.100 61.800 26.200 ;
        RECT 63.800 26.100 64.100 26.800 ;
        RECT 61.400 25.800 64.100 26.100 ;
        RECT 65.400 26.100 65.800 26.200 ;
        RECT 71.000 26.100 71.400 26.200 ;
        RECT 65.400 25.800 71.400 26.100 ;
        RECT 84.600 26.100 85.000 26.200 ;
        RECT 94.200 26.100 94.600 26.200 ;
        RECT 84.600 25.800 94.600 26.100 ;
        RECT 95.000 26.100 95.400 26.200 ;
        RECT 96.600 26.100 97.000 26.200 ;
        RECT 95.000 25.800 97.000 26.100 ;
        RECT 50.200 25.200 50.500 25.800 ;
        RECT 8.600 24.800 9.000 25.200 ;
        RECT 15.000 24.800 15.400 25.200 ;
        RECT 15.800 25.100 16.200 25.200 ;
        RECT 20.600 25.100 21.000 25.200 ;
        RECT 15.800 24.800 21.000 25.100 ;
        RECT 27.800 25.100 28.200 25.200 ;
        RECT 32.600 25.100 33.000 25.200 ;
        RECT 35.800 25.100 36.200 25.200 ;
        RECT 27.800 24.800 36.200 25.100 ;
        RECT 38.200 25.100 38.600 25.200 ;
        RECT 43.000 25.100 43.400 25.200 ;
        RECT 38.200 24.800 43.400 25.100 ;
        RECT 50.200 24.800 50.600 25.200 ;
        RECT 51.000 25.100 51.400 25.200 ;
        RECT 53.400 25.100 53.800 25.200 ;
        RECT 51.000 24.800 53.800 25.100 ;
        RECT 54.200 25.100 54.600 25.200 ;
        RECT 69.400 25.100 69.800 25.200 ;
        RECT 54.200 24.800 69.800 25.100 ;
        RECT 87.000 25.100 87.400 25.200 ;
        RECT 88.600 25.100 89.000 25.200 ;
        RECT 95.800 25.100 96.200 25.200 ;
        RECT 87.000 24.800 96.200 25.100 ;
        RECT 8.600 24.200 8.900 24.800 ;
        RECT 15.000 24.200 15.300 24.800 ;
        RECT 3.000 24.100 3.400 24.200 ;
        RECT 5.400 24.100 5.800 24.200 ;
        RECT 3.000 23.800 5.800 24.100 ;
        RECT 8.600 23.800 9.000 24.200 ;
        RECT 15.000 23.800 15.400 24.200 ;
        RECT 15.800 24.100 16.200 24.200 ;
        RECT 27.800 24.100 28.200 24.200 ;
        RECT 15.800 23.800 28.200 24.100 ;
        RECT 39.000 24.100 39.400 24.200 ;
        RECT 49.400 24.100 49.800 24.200 ;
        RECT 50.200 24.100 50.600 24.200 ;
        RECT 39.000 23.800 50.600 24.100 ;
        RECT 56.600 24.100 57.000 24.200 ;
        RECT 75.000 24.100 75.400 24.200 ;
        RECT 79.000 24.100 79.400 24.200 ;
        RECT 79.800 24.100 80.200 24.200 ;
        RECT 56.600 23.800 88.100 24.100 ;
        RECT 87.800 23.200 88.100 23.800 ;
        RECT 7.000 22.800 7.400 23.200 ;
        RECT 23.800 23.100 24.200 23.200 ;
        RECT 33.400 23.100 33.800 23.200 ;
        RECT 23.000 22.800 33.800 23.100 ;
        RECT 47.800 23.100 48.200 23.200 ;
        RECT 50.200 23.100 50.600 23.200 ;
        RECT 47.800 22.800 50.600 23.100 ;
        RECT 75.000 23.100 75.400 23.200 ;
        RECT 83.000 23.100 83.400 23.200 ;
        RECT 75.000 22.800 83.400 23.100 ;
        RECT 87.800 22.800 88.200 23.200 ;
        RECT 7.000 22.100 7.300 22.800 ;
        RECT 43.000 22.100 43.400 22.200 ;
        RECT 7.000 21.800 43.400 22.100 ;
        RECT 43.800 22.100 44.200 22.200 ;
        RECT 58.200 22.100 58.600 22.200 ;
        RECT 43.800 21.800 58.600 22.100 ;
        RECT 34.200 21.100 34.600 21.200 ;
        RECT 54.200 21.100 54.600 21.200 ;
        RECT 34.200 20.800 54.600 21.100 ;
        RECT 36.600 20.100 37.000 20.200 ;
        RECT 65.400 20.100 65.800 20.200 ;
        RECT 66.200 20.100 66.600 20.200 ;
        RECT 36.600 19.800 66.600 20.100 ;
        RECT 9.400 19.100 9.800 19.200 ;
        RECT 31.800 19.100 32.200 19.200 ;
        RECT 9.400 18.800 32.200 19.100 ;
        RECT 32.600 19.100 33.000 19.200 ;
        RECT 43.000 19.100 43.400 19.200 ;
        RECT 57.400 19.100 57.800 19.200 ;
        RECT 32.600 18.800 57.800 19.100 ;
        RECT 61.400 18.800 61.800 19.200 ;
        RECT 23.000 17.800 23.400 18.200 ;
        RECT 61.400 18.100 61.700 18.800 ;
        RECT 91.000 18.100 91.400 18.200 ;
        RECT 61.400 17.800 91.400 18.100 ;
        RECT 23.000 17.200 23.300 17.800 ;
        RECT 7.800 16.800 11.300 17.100 ;
        RECT 7.800 16.200 8.100 16.800 ;
        RECT 11.000 16.200 11.300 16.800 ;
        RECT 12.600 16.800 13.000 17.200 ;
        RECT 19.000 17.100 19.400 17.200 ;
        RECT 23.000 17.100 23.400 17.200 ;
        RECT 30.200 17.100 30.600 17.200 ;
        RECT 19.000 16.800 30.600 17.100 ;
        RECT 33.400 17.100 33.800 17.200 ;
        RECT 38.200 17.100 38.600 17.200 ;
        RECT 33.400 16.800 38.600 17.100 ;
        RECT 48.600 16.800 49.000 17.200 ;
        RECT 50.200 16.800 50.600 17.200 ;
        RECT 84.600 16.800 85.000 17.200 ;
        RECT 7.800 15.800 8.200 16.200 ;
        RECT 11.000 15.800 11.400 16.200 ;
        RECT 12.600 16.100 12.900 16.800 ;
        RECT 15.000 16.100 15.400 16.200 ;
        RECT 12.600 15.800 15.400 16.100 ;
        RECT 18.200 16.100 18.600 16.200 ;
        RECT 19.000 16.100 19.400 16.200 ;
        RECT 18.200 15.800 19.400 16.100 ;
        RECT 21.400 16.100 21.800 16.200 ;
        RECT 22.200 16.100 22.600 16.200 ;
        RECT 35.800 16.100 36.200 16.200 ;
        RECT 21.400 15.800 36.200 16.100 ;
        RECT 48.600 16.100 48.900 16.800 ;
        RECT 50.200 16.100 50.500 16.800 ;
        RECT 84.600 16.200 84.900 16.800 ;
        RECT 48.600 15.800 50.500 16.100 ;
        RECT 59.000 15.800 59.400 16.200 ;
        RECT 63.000 16.100 63.400 16.200 ;
        RECT 79.000 16.100 79.400 16.200 ;
        RECT 63.000 15.800 79.400 16.100 ;
        RECT 82.200 16.100 82.600 16.200 ;
        RECT 83.800 16.100 84.200 16.200 ;
        RECT 82.200 15.800 84.200 16.100 ;
        RECT 84.600 15.800 85.000 16.200 ;
        RECT 92.600 16.100 93.000 16.200 ;
        RECT 94.200 16.100 94.600 16.200 ;
        RECT 92.600 15.800 94.600 16.100 ;
        RECT 59.000 15.200 59.300 15.800 ;
        RECT 12.600 15.100 13.000 15.200 ;
        RECT 13.400 15.100 13.800 15.200 ;
        RECT 12.600 14.800 13.800 15.100 ;
        RECT 15.800 15.100 16.200 15.200 ;
        RECT 49.400 15.100 49.800 15.200 ;
        RECT 51.800 15.100 52.200 15.200 ;
        RECT 15.800 14.800 52.200 15.100 ;
        RECT 59.000 14.800 59.400 15.200 ;
        RECT 63.000 15.100 63.400 15.200 ;
        RECT 75.800 15.100 76.200 15.200 ;
        RECT 63.000 14.800 76.200 15.100 ;
        RECT 79.000 15.100 79.400 15.200 ;
        RECT 82.200 15.100 82.600 15.200 ;
        RECT 79.000 14.800 82.600 15.100 ;
        RECT 83.000 15.100 83.400 15.200 ;
        RECT 87.800 15.100 88.200 15.200 ;
        RECT 88.600 15.100 89.000 15.200 ;
        RECT 83.000 14.800 89.000 15.100 ;
        RECT 91.000 15.100 91.400 15.200 ;
        RECT 92.600 15.100 93.000 15.200 ;
        RECT 91.000 14.800 93.000 15.100 ;
        RECT 4.600 14.100 5.000 14.200 ;
        RECT 5.400 14.100 5.800 14.200 ;
        RECT 4.600 13.800 5.800 14.100 ;
        RECT 30.200 14.100 30.600 14.200 ;
        RECT 42.200 14.100 42.600 14.200 ;
        RECT 30.200 13.800 42.600 14.100 ;
        RECT 43.000 14.100 43.400 14.200 ;
        RECT 47.000 14.100 47.400 14.200 ;
        RECT 43.000 13.800 47.400 14.100 ;
        RECT 57.400 14.100 57.800 14.200 ;
        RECT 62.200 14.100 62.600 14.200 ;
        RECT 57.400 13.800 62.600 14.100 ;
        RECT 63.800 14.100 64.200 14.200 ;
        RECT 71.800 14.100 72.200 14.200 ;
        RECT 76.600 14.100 77.000 14.200 ;
        RECT 78.200 14.100 78.600 14.200 ;
        RECT 83.800 14.100 84.200 14.200 ;
        RECT 87.000 14.100 87.400 14.200 ;
        RECT 63.800 13.800 87.400 14.100 ;
        RECT 4.600 13.100 5.000 13.200 ;
        RECT 9.400 13.100 9.800 13.200 ;
        RECT 4.600 12.800 9.800 13.100 ;
        RECT 10.200 13.100 10.600 13.200 ;
        RECT 12.600 13.100 13.000 13.200 ;
        RECT 10.200 12.800 13.000 13.100 ;
        RECT 13.400 13.100 13.800 13.200 ;
        RECT 24.600 13.100 25.000 13.200 ;
        RECT 25.400 13.100 25.800 13.200 ;
        RECT 13.400 12.800 20.100 13.100 ;
        RECT 24.600 12.800 25.800 13.100 ;
        RECT 36.600 12.800 37.000 13.200 ;
        RECT 39.000 13.100 39.400 13.200 ;
        RECT 41.400 13.100 41.800 13.200 ;
        RECT 39.000 12.800 41.800 13.100 ;
        RECT 42.200 13.100 42.500 13.800 ;
        RECT 53.400 13.100 53.800 13.200 ;
        RECT 67.800 13.100 68.200 13.200 ;
        RECT 42.200 12.800 53.800 13.100 ;
        RECT 65.400 12.800 68.200 13.100 ;
        RECT 68.600 13.100 69.000 13.200 ;
        RECT 73.400 13.100 73.800 13.200 ;
        RECT 68.600 12.800 73.800 13.100 ;
        RECT 76.600 13.100 77.000 13.200 ;
        RECT 80.600 13.100 81.000 13.200 ;
        RECT 76.600 12.800 81.000 13.100 ;
        RECT 82.200 13.100 82.600 13.200 ;
        RECT 83.000 13.100 83.400 13.200 ;
        RECT 82.200 12.800 83.400 13.100 ;
        RECT 85.400 13.100 85.800 13.200 ;
        RECT 89.400 13.100 89.800 13.200 ;
        RECT 90.200 13.100 90.600 13.200 ;
        RECT 85.400 12.800 90.600 13.100 ;
        RECT 19.800 12.200 20.100 12.800 ;
        RECT 16.600 12.100 17.000 12.200 ;
        RECT 19.000 12.100 19.400 12.200 ;
        RECT 16.600 11.800 19.400 12.100 ;
        RECT 19.800 11.800 20.200 12.200 ;
        RECT 36.600 12.100 36.900 12.800 ;
        RECT 65.400 12.200 65.700 12.800 ;
        RECT 39.800 12.100 40.200 12.200 ;
        RECT 41.400 12.100 41.800 12.200 ;
        RECT 43.800 12.100 44.200 12.200 ;
        RECT 36.600 11.800 40.200 12.100 ;
        RECT 40.600 11.800 44.200 12.100 ;
        RECT 45.400 12.100 45.800 12.200 ;
        RECT 56.600 12.100 57.000 12.200 ;
        RECT 45.400 11.800 57.000 12.100 ;
        RECT 65.400 11.800 65.800 12.200 ;
        RECT 67.000 12.100 67.400 12.200 ;
        RECT 74.200 12.100 74.600 12.200 ;
        RECT 66.200 11.800 74.600 12.100 ;
        RECT 75.000 12.100 75.400 12.200 ;
        RECT 77.400 12.100 77.800 12.200 ;
        RECT 80.600 12.100 81.000 12.200 ;
        RECT 92.600 12.100 93.000 12.200 ;
        RECT 75.000 11.800 77.800 12.100 ;
        RECT 79.800 11.800 93.000 12.100 ;
        RECT 3.800 11.100 4.200 11.200 ;
        RECT 18.200 11.100 18.600 11.200 ;
        RECT 23.800 11.100 24.200 11.200 ;
        RECT 28.600 11.100 29.000 11.200 ;
        RECT 31.000 11.100 31.400 11.200 ;
        RECT 3.800 10.800 31.400 11.100 ;
        RECT 31.800 11.100 32.200 11.200 ;
        RECT 40.600 11.100 41.000 11.200 ;
        RECT 67.000 11.100 67.400 11.200 ;
        RECT 31.800 10.800 67.400 11.100 ;
        RECT 8.600 10.100 9.000 10.200 ;
        RECT 13.400 10.100 13.800 10.200 ;
        RECT 8.600 9.800 13.800 10.100 ;
        RECT 15.800 10.100 16.200 10.200 ;
        RECT 26.200 10.100 26.600 10.200 ;
        RECT 32.600 10.100 33.000 10.200 ;
        RECT 34.200 10.100 34.600 10.200 ;
        RECT 15.800 9.800 34.600 10.100 ;
        RECT 50.200 9.800 50.600 10.200 ;
        RECT 53.400 10.100 53.800 10.200 ;
        RECT 58.200 10.100 58.600 10.200 ;
        RECT 53.400 9.800 58.600 10.100 ;
        RECT 13.400 9.100 13.700 9.800 ;
        RECT 50.200 9.200 50.500 9.800 ;
        RECT 23.800 9.100 24.200 9.200 ;
        RECT 37.400 9.100 37.800 9.200 ;
        RECT 13.400 8.800 37.800 9.100 ;
        RECT 38.200 9.100 38.600 9.200 ;
        RECT 45.400 9.100 45.800 9.200 ;
        RECT 38.200 8.800 45.800 9.100 ;
        RECT 50.200 8.800 50.600 9.200 ;
        RECT 61.400 9.100 61.800 9.200 ;
        RECT 63.800 9.100 64.200 9.200 ;
        RECT 61.400 8.800 64.200 9.100 ;
        RECT 64.600 9.100 65.000 9.200 ;
        RECT 76.600 9.100 77.000 9.200 ;
        RECT 64.600 8.800 77.000 9.100 ;
        RECT 84.600 9.100 85.000 9.200 ;
        RECT 95.000 9.100 95.400 9.200 ;
        RECT 84.600 8.800 95.400 9.100 ;
        RECT 55.000 8.100 55.400 8.200 ;
        RECT 69.400 8.100 69.800 8.200 ;
        RECT 78.200 8.100 78.600 8.200 ;
        RECT 55.000 7.800 78.600 8.100 ;
        RECT 27.000 7.100 27.400 7.200 ;
        RECT 27.800 7.100 28.200 7.200 ;
        RECT 27.000 6.800 28.200 7.100 ;
        RECT 43.800 7.100 44.200 7.200 ;
        RECT 44.600 7.100 45.000 7.200 ;
        RECT 63.800 7.100 64.200 7.200 ;
        RECT 43.800 6.800 64.200 7.100 ;
        RECT 74.200 7.100 74.600 7.200 ;
        RECT 84.600 7.100 85.000 7.200 ;
        RECT 74.200 6.800 85.000 7.100 ;
        RECT 12.600 6.100 13.000 6.200 ;
        RECT 14.200 6.100 14.600 6.200 ;
        RECT 12.600 5.800 14.600 6.100 ;
        RECT 27.000 6.100 27.400 6.200 ;
        RECT 30.200 6.100 30.600 6.200 ;
        RECT 27.000 5.800 30.600 6.100 ;
        RECT 34.200 5.800 34.600 6.200 ;
        RECT 64.600 6.100 65.000 6.200 ;
        RECT 65.400 6.100 65.800 6.200 ;
        RECT 77.400 6.100 77.800 6.200 ;
        RECT 64.600 5.800 65.800 6.100 ;
        RECT 72.600 5.800 77.800 6.100 ;
        RECT 79.000 6.100 79.400 6.200 ;
        RECT 79.000 5.800 80.900 6.100 ;
        RECT 18.200 5.100 18.600 5.200 ;
        RECT 20.600 5.100 21.000 5.200 ;
        RECT 34.200 5.100 34.500 5.800 ;
        RECT 72.600 5.200 72.900 5.800 ;
        RECT 80.600 5.200 80.900 5.800 ;
        RECT 18.200 4.800 34.500 5.100 ;
        RECT 37.400 5.100 37.800 5.200 ;
        RECT 41.400 5.100 41.800 5.200 ;
        RECT 37.400 4.800 41.800 5.100 ;
        RECT 72.600 4.800 73.000 5.200 ;
        RECT 79.000 5.100 79.400 5.200 ;
        RECT 79.800 5.100 80.200 5.200 ;
        RECT 79.000 4.800 80.200 5.100 ;
        RECT 80.600 4.800 81.000 5.200 ;
        RECT 19.000 4.100 19.400 4.200 ;
        RECT 36.600 4.100 37.000 4.200 ;
        RECT 19.000 3.800 37.000 4.100 ;
        RECT 77.400 4.100 77.800 4.200 ;
        RECT 83.800 4.100 84.200 4.200 ;
        RECT 77.400 3.800 84.200 4.100 ;
      LAYER via3 ;
        RECT 75.800 76.800 76.200 77.200 ;
        RECT 70.200 72.800 70.600 73.200 ;
        RECT 61.400 71.800 61.800 72.200 ;
        RECT 47.000 70.800 47.400 71.200 ;
        RECT 70.200 67.800 70.600 68.200 ;
        RECT 66.200 66.800 66.600 67.200 ;
        RECT 43.800 65.800 44.200 66.200 ;
        RECT 79.000 61.800 79.400 62.200 ;
        RECT 84.600 61.800 85.000 62.200 ;
        RECT 47.800 60.800 48.200 61.200 ;
        RECT 61.400 58.800 61.800 59.200 ;
        RECT 95.800 54.800 96.200 55.200 ;
        RECT 51.800 52.800 52.200 53.200 ;
        RECT 64.600 52.800 65.000 53.200 ;
        RECT 62.200 51.800 62.600 52.200 ;
        RECT 11.000 50.800 11.400 51.200 ;
        RECT 51.000 50.800 51.400 51.200 ;
        RECT 45.400 49.800 45.800 50.200 ;
        RECT 54.200 49.800 54.600 50.200 ;
        RECT 67.000 49.800 67.400 50.200 ;
        RECT 83.800 47.800 84.200 48.200 ;
        RECT 63.000 46.800 63.400 47.200 ;
        RECT 81.400 46.800 81.800 47.200 ;
        RECT 81.400 45.800 81.800 46.200 ;
        RECT 7.800 43.800 8.200 44.200 ;
        RECT 3.800 40.800 4.200 41.200 ;
        RECT 23.000 37.800 23.400 38.200 ;
        RECT 95.000 37.800 95.400 38.200 ;
        RECT 14.200 34.800 14.600 35.200 ;
        RECT 50.200 34.800 50.600 35.200 ;
        RECT 70.200 33.800 70.600 34.200 ;
        RECT 24.600 32.800 25.000 33.200 ;
        RECT 41.400 32.800 41.800 33.200 ;
        RECT 19.000 30.800 19.400 31.200 ;
        RECT 62.200 29.800 62.600 30.200 ;
        RECT 43.000 28.800 43.400 29.200 ;
        RECT 59.800 28.800 60.200 29.200 ;
        RECT 63.000 28.800 63.400 29.200 ;
        RECT 42.200 27.800 42.600 28.200 ;
        RECT 19.800 26.800 20.200 27.200 ;
        RECT 23.800 26.800 24.200 27.200 ;
        RECT 38.200 26.800 38.600 27.200 ;
        RECT 60.600 26.800 61.000 27.200 ;
        RECT 62.200 26.800 62.600 27.200 ;
        RECT 59.800 25.800 60.200 26.200 ;
        RECT 53.400 24.800 53.800 25.200 ;
        RECT 95.800 24.800 96.200 25.200 ;
        RECT 50.200 23.800 50.600 24.200 ;
        RECT 79.800 23.800 80.200 24.200 ;
        RECT 83.000 22.800 83.400 23.200 ;
        RECT 43.000 21.800 43.400 22.200 ;
        RECT 66.200 19.800 66.600 20.200 ;
        RECT 31.800 18.800 32.200 19.200 ;
        RECT 19.000 15.800 19.400 16.200 ;
        RECT 22.200 15.800 22.600 16.200 ;
        RECT 49.400 14.800 49.800 15.200 ;
        RECT 88.600 14.800 89.000 15.200 ;
        RECT 83.000 12.800 83.400 13.200 ;
        RECT 90.200 12.800 90.600 13.200 ;
        RECT 74.200 11.800 74.600 12.200 ;
        RECT 18.200 10.800 18.600 11.200 ;
        RECT 67.000 10.800 67.400 11.200 ;
        RECT 95.000 8.800 95.400 9.200 ;
        RECT 65.400 5.800 65.800 6.200 ;
        RECT 79.800 4.800 80.200 5.200 ;
      LAYER metal4 ;
        RECT 75.800 76.800 76.200 77.200 ;
        RECT 61.400 72.800 61.800 73.200 ;
        RECT 62.200 72.800 62.600 73.200 ;
        RECT 70.200 72.800 70.600 73.200 ;
        RECT 61.400 72.200 61.700 72.800 ;
        RECT 61.400 71.800 61.800 72.200 ;
        RECT 3.800 70.800 4.200 71.200 ;
        RECT 47.000 70.800 47.400 71.200 ;
        RECT 3.800 41.200 4.100 70.800 ;
        RECT 4.600 68.800 5.000 69.200 ;
        RECT 3.800 40.800 4.200 41.200 ;
        RECT 4.600 30.200 4.900 68.800 ;
        RECT 43.800 65.800 44.200 66.200 ;
        RECT 7.000 64.800 7.400 65.200 ;
        RECT 15.000 64.800 15.400 65.200 ;
        RECT 7.000 59.200 7.300 64.800 ;
        RECT 7.800 60.800 8.200 61.200 ;
        RECT 7.000 58.800 7.400 59.200 ;
        RECT 7.000 42.200 7.300 58.800 ;
        RECT 7.800 44.200 8.100 60.800 ;
        RECT 11.000 51.100 11.400 51.200 ;
        RECT 10.200 50.800 11.400 51.100 ;
        RECT 7.800 43.800 8.200 44.200 ;
        RECT 7.000 41.800 7.400 42.200 ;
        RECT 4.600 29.800 5.000 30.200 ;
        RECT 7.800 26.200 8.100 43.800 ;
        RECT 10.200 37.200 10.500 50.800 ;
        RECT 10.200 36.800 10.600 37.200 ;
        RECT 14.200 34.800 14.600 35.200 ;
        RECT 14.200 27.200 14.500 34.800 ;
        RECT 14.200 26.800 14.600 27.200 ;
        RECT 7.800 25.800 8.200 26.200 ;
        RECT 15.000 25.200 15.300 64.800 ;
        RECT 22.200 63.800 22.600 64.200 ;
        RECT 22.200 57.200 22.500 63.800 ;
        RECT 22.200 56.800 22.600 57.200 ;
        RECT 19.000 30.800 19.400 31.200 ;
        RECT 8.600 25.100 9.000 25.200 ;
        RECT 9.400 25.100 9.800 25.200 ;
        RECT 8.600 24.800 9.800 25.100 ;
        RECT 15.000 24.800 15.400 25.200 ;
        RECT 15.800 24.800 16.200 25.200 ;
        RECT 15.800 24.200 16.100 24.800 ;
        RECT 15.800 23.800 16.200 24.200 ;
        RECT 19.000 16.200 19.300 30.800 ;
        RECT 19.800 27.100 20.200 27.200 ;
        RECT 20.600 27.100 21.000 27.200 ;
        RECT 19.800 26.800 21.000 27.100 ;
        RECT 22.200 16.200 22.500 56.800 ;
        RECT 43.800 48.200 44.100 65.800 ;
        RECT 45.400 49.800 45.800 50.200 ;
        RECT 43.800 47.800 44.200 48.200 ;
        RECT 38.200 46.800 38.600 47.200 ;
        RECT 38.200 44.200 38.500 46.800 ;
        RECT 38.200 43.800 38.600 44.200 ;
        RECT 23.000 37.800 23.400 38.200 ;
        RECT 23.800 37.800 24.200 38.200 ;
        RECT 23.000 18.200 23.300 37.800 ;
        RECT 23.800 27.200 24.100 37.800 ;
        RECT 43.000 35.800 43.400 36.200 ;
        RECT 24.600 32.800 25.000 33.200 ;
        RECT 41.400 33.100 41.800 33.200 ;
        RECT 42.200 33.100 42.600 33.200 ;
        RECT 41.400 32.800 42.600 33.100 ;
        RECT 23.800 26.800 24.200 27.200 ;
        RECT 23.000 17.800 23.400 18.200 ;
        RECT 19.000 16.100 19.400 16.200 ;
        RECT 18.200 15.800 19.400 16.100 ;
        RECT 22.200 15.800 22.600 16.200 ;
        RECT 4.600 14.100 5.000 14.200 ;
        RECT 5.400 14.100 5.800 14.200 ;
        RECT 4.600 13.800 5.800 14.100 ;
        RECT 13.400 13.800 13.800 14.200 ;
        RECT 13.400 13.200 13.700 13.800 ;
        RECT 13.400 12.800 13.800 13.200 ;
        RECT 18.200 11.200 18.500 15.800 ;
        RECT 24.600 13.200 24.900 32.800 ;
        RECT 43.000 29.200 43.300 35.800 ;
        RECT 43.000 28.800 43.400 29.200 ;
        RECT 43.000 28.200 43.300 28.800 ;
        RECT 42.200 27.800 42.600 28.200 ;
        RECT 43.000 27.800 43.400 28.200 ;
        RECT 38.200 26.800 38.600 27.200 ;
        RECT 38.200 25.200 38.500 26.800 ;
        RECT 42.200 26.200 42.500 27.800 ;
        RECT 42.200 25.800 42.600 26.200 ;
        RECT 38.200 24.800 38.600 25.200 ;
        RECT 43.000 21.800 43.400 22.200 ;
        RECT 31.800 18.800 32.200 19.200 ;
        RECT 24.600 12.800 25.000 13.200 ;
        RECT 31.800 11.200 32.100 18.800 ;
        RECT 43.000 15.200 43.300 21.800 ;
        RECT 43.000 14.800 43.400 15.200 ;
        RECT 18.200 10.800 18.600 11.200 ;
        RECT 31.800 10.800 32.200 11.200 ;
        RECT 38.200 8.800 38.600 9.200 ;
        RECT 38.200 7.200 38.500 8.800 ;
        RECT 43.800 7.200 44.100 47.800 ;
        RECT 44.600 32.800 45.000 33.200 ;
        RECT 44.600 28.200 44.900 32.800 ;
        RECT 44.600 27.800 45.000 28.200 ;
        RECT 45.400 12.200 45.700 49.800 ;
        RECT 47.000 37.200 47.300 70.800 ;
        RECT 51.000 61.800 51.400 62.200 ;
        RECT 47.800 60.800 48.200 61.200 ;
        RECT 47.000 36.800 47.400 37.200 ;
        RECT 47.800 26.200 48.100 60.800 ;
        RECT 51.000 51.200 51.300 61.800 ;
        RECT 61.400 58.800 61.800 59.200 ;
        RECT 51.800 52.800 52.200 53.200 ;
        RECT 51.000 50.800 51.400 51.200 ;
        RECT 51.800 45.200 52.100 52.800 ;
        RECT 54.200 50.100 54.600 50.200 ;
        RECT 53.400 49.800 54.600 50.100 ;
        RECT 53.400 45.200 53.700 49.800 ;
        RECT 51.800 44.800 52.200 45.200 ;
        RECT 53.400 44.800 53.800 45.200 ;
        RECT 53.400 37.800 53.800 38.200 ;
        RECT 50.200 35.100 50.600 35.200 ;
        RECT 49.400 34.800 50.600 35.100 ;
        RECT 47.800 25.800 48.200 26.200 ;
        RECT 49.400 15.200 49.700 34.800 ;
        RECT 53.400 25.200 53.700 37.800 ;
        RECT 56.600 28.800 57.000 29.200 ;
        RECT 59.800 29.100 60.200 29.200 ;
        RECT 60.600 29.100 61.000 29.200 ;
        RECT 59.800 28.800 61.000 29.100 ;
        RECT 53.400 24.800 53.800 25.200 ;
        RECT 56.600 24.200 56.900 28.800 ;
        RECT 59.800 27.100 60.200 27.200 ;
        RECT 60.600 27.100 61.000 27.200 ;
        RECT 59.800 26.800 61.000 27.100 ;
        RECT 61.400 26.200 61.700 58.800 ;
        RECT 62.200 52.200 62.500 72.800 ;
        RECT 70.200 68.200 70.500 72.800 ;
        RECT 70.200 67.800 70.600 68.200 ;
        RECT 66.200 66.800 66.600 67.200 ;
        RECT 64.600 53.100 65.000 53.200 ;
        RECT 63.800 52.800 65.000 53.100 ;
        RECT 62.200 51.800 62.600 52.200 ;
        RECT 63.000 47.100 63.400 47.200 ;
        RECT 63.800 47.100 64.100 52.800 ;
        RECT 63.000 46.800 64.100 47.100 ;
        RECT 62.200 46.100 62.600 46.200 ;
        RECT 62.200 45.800 63.300 46.100 ;
        RECT 62.200 29.800 62.600 30.200 ;
        RECT 62.200 27.200 62.500 29.800 ;
        RECT 63.000 29.200 63.300 45.800 ;
        RECT 63.800 39.200 64.100 46.800 ;
        RECT 63.800 38.800 64.200 39.200 ;
        RECT 63.000 28.800 63.400 29.200 ;
        RECT 62.200 26.800 62.600 27.200 ;
        RECT 59.000 26.100 59.400 26.200 ;
        RECT 59.800 26.100 60.200 26.200 ;
        RECT 59.000 25.800 60.200 26.100 ;
        RECT 61.400 25.800 61.800 26.200 ;
        RECT 50.200 23.800 50.600 24.200 ;
        RECT 56.600 23.800 57.000 24.200 ;
        RECT 49.400 14.800 49.800 15.200 ;
        RECT 45.400 11.800 45.800 12.200 ;
        RECT 50.200 9.200 50.500 23.800 ;
        RECT 66.200 20.200 66.500 66.800 ;
        RECT 67.000 49.800 67.400 50.200 ;
        RECT 67.000 48.200 67.300 49.800 ;
        RECT 67.000 47.800 67.400 48.200 ;
        RECT 75.800 42.200 76.100 76.800 ;
        RECT 79.000 73.800 79.400 74.200 ;
        RECT 79.000 62.200 79.300 73.800 ;
        RECT 81.400 73.100 81.800 73.200 ;
        RECT 82.200 73.100 82.600 73.200 ;
        RECT 81.400 72.800 82.600 73.100 ;
        RECT 79.000 61.800 79.400 62.200 ;
        RECT 84.600 61.800 85.000 62.200 ;
        RECT 90.200 61.800 90.600 62.200 ;
        RECT 83.800 47.800 84.200 48.200 ;
        RECT 80.600 47.100 81.000 47.200 ;
        RECT 81.400 47.100 81.800 47.200 ;
        RECT 80.600 46.800 81.800 47.100 ;
        RECT 82.200 46.800 82.600 47.200 ;
        RECT 81.400 46.100 81.800 46.200 ;
        RECT 82.200 46.100 82.500 46.800 ;
        RECT 81.400 45.800 82.500 46.100 ;
        RECT 75.800 41.800 76.200 42.200 ;
        RECT 67.000 35.800 67.400 36.200 ;
        RECT 66.200 19.800 66.600 20.200 ;
        RECT 58.200 15.100 58.600 15.200 ;
        RECT 59.000 15.100 59.400 15.200 ;
        RECT 58.200 14.800 59.400 15.100 ;
        RECT 67.000 11.200 67.300 35.800 ;
        RECT 83.000 35.100 83.400 35.200 ;
        RECT 83.800 35.100 84.100 47.800 ;
        RECT 83.000 34.800 84.100 35.100 ;
        RECT 70.200 33.800 70.600 34.200 ;
        RECT 70.200 30.200 70.500 33.800 ;
        RECT 82.200 33.100 82.600 33.200 ;
        RECT 82.200 32.800 83.300 33.100 ;
        RECT 72.600 30.800 73.000 31.200 ;
        RECT 70.200 29.800 70.600 30.200 ;
        RECT 72.600 29.200 72.900 30.800 ;
        RECT 72.600 28.800 73.000 29.200 ;
        RECT 79.800 23.800 80.200 24.200 ;
        RECT 74.200 11.800 74.600 12.200 ;
        RECT 67.000 10.800 67.400 11.200 ;
        RECT 50.200 8.800 50.600 9.200 ;
        RECT 64.600 8.800 65.000 9.200 ;
        RECT 27.000 7.100 27.400 7.200 ;
        RECT 27.800 7.100 28.200 7.200 ;
        RECT 27.000 6.800 28.200 7.100 ;
        RECT 38.200 6.800 38.600 7.200 ;
        RECT 43.800 6.800 44.200 7.200 ;
        RECT 64.600 6.100 64.900 8.800 ;
        RECT 74.200 7.200 74.500 11.800 ;
        RECT 74.200 6.800 74.600 7.200 ;
        RECT 65.400 6.100 65.800 6.200 ;
        RECT 64.600 5.800 65.800 6.100 ;
        RECT 79.800 5.200 80.100 23.800 ;
        RECT 83.000 23.200 83.300 32.800 ;
        RECT 84.600 26.200 84.900 61.800 ;
        RECT 88.600 47.800 89.000 48.200 ;
        RECT 84.600 25.800 85.000 26.200 ;
        RECT 83.000 22.800 83.400 23.200 ;
        RECT 84.600 17.200 84.900 25.800 ;
        RECT 84.600 16.800 85.000 17.200 ;
        RECT 82.200 15.800 82.600 16.200 ;
        RECT 82.200 13.100 82.500 15.800 ;
        RECT 88.600 15.200 88.900 47.800 ;
        RECT 89.400 45.800 89.800 46.200 ;
        RECT 89.400 33.200 89.700 45.800 ;
        RECT 89.400 32.800 89.800 33.200 ;
        RECT 88.600 14.800 89.000 15.200 ;
        RECT 90.200 13.200 90.500 61.800 ;
        RECT 95.800 54.800 96.200 55.200 ;
        RECT 95.000 37.800 95.400 38.200 ;
        RECT 95.000 26.200 95.300 37.800 ;
        RECT 95.000 25.800 95.400 26.200 ;
        RECT 83.000 13.100 83.400 13.200 ;
        RECT 82.200 12.800 83.400 13.100 ;
        RECT 90.200 12.800 90.600 13.200 ;
        RECT 95.000 9.200 95.300 25.800 ;
        RECT 95.800 25.200 96.100 54.800 ;
        RECT 95.800 24.800 96.200 25.200 ;
        RECT 95.000 8.800 95.400 9.200 ;
        RECT 79.800 4.800 80.200 5.200 ;
      LAYER via4 ;
        RECT 9.400 24.800 9.800 25.200 ;
        RECT 20.600 26.800 21.000 27.200 ;
        RECT 42.200 32.800 42.600 33.200 ;
        RECT 5.400 13.800 5.800 14.200 ;
        RECT 60.600 28.800 61.000 29.200 ;
        RECT 27.800 6.800 28.200 7.200 ;
      LAYER metal5 ;
        RECT 61.400 73.100 61.800 73.200 ;
        RECT 81.400 73.100 81.800 73.200 ;
        RECT 61.400 72.800 81.800 73.100 ;
        RECT 38.200 47.100 38.600 47.200 ;
        RECT 80.600 47.100 81.000 47.200 ;
        RECT 38.200 46.800 81.000 47.100 ;
        RECT 42.200 33.100 42.600 33.200 ;
        RECT 44.600 33.100 45.000 33.200 ;
        RECT 42.200 32.800 45.000 33.100 ;
        RECT 60.600 29.100 61.000 29.200 ;
        RECT 72.600 29.100 73.000 29.200 ;
        RECT 60.600 28.800 73.000 29.100 ;
        RECT 20.600 27.100 21.000 27.200 ;
        RECT 59.800 27.100 60.200 27.200 ;
        RECT 20.600 26.800 60.200 27.100 ;
        RECT 42.200 26.100 42.600 26.200 ;
        RECT 59.000 26.100 59.400 26.200 ;
        RECT 42.200 25.800 59.400 26.100 ;
        RECT 9.400 25.100 9.800 25.200 ;
        RECT 15.800 25.100 16.200 25.200 ;
        RECT 9.400 24.800 16.200 25.100 ;
        RECT 43.000 15.100 43.400 15.200 ;
        RECT 58.200 15.100 58.600 15.200 ;
        RECT 43.000 14.800 58.600 15.100 ;
        RECT 5.400 14.100 5.800 14.200 ;
        RECT 13.400 14.100 13.800 14.200 ;
        RECT 5.400 13.800 13.800 14.100 ;
        RECT 27.800 7.100 28.200 7.200 ;
        RECT 38.200 7.100 38.600 7.200 ;
        RECT 27.800 6.800 38.600 7.100 ;
  END
END ALU
END LIBRARY

