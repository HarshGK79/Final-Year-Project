magic
tech scmos
timestamp 1744883066
<< metal1 >>
rect 272 803 274 807
rect 278 803 281 807
rect 285 803 288 807
rect 133 768 134 772
rect 102 766 106 768
rect 54 758 65 761
rect 102 758 110 761
rect 214 758 225 761
rect 274 758 297 761
rect 22 748 33 751
rect 246 748 254 751
rect 366 751 370 754
rect 362 748 370 751
rect 430 748 446 751
rect 462 748 473 751
rect 590 748 614 751
rect 734 748 742 751
rect 774 751 778 754
rect 774 748 782 751
rect 852 748 881 751
rect 246 746 250 748
rect 142 738 150 741
rect 182 738 201 741
rect 318 738 337 741
rect 414 738 433 741
rect 518 738 534 741
rect 542 738 550 741
rect 606 738 633 741
rect 638 738 657 741
rect 798 738 833 741
rect 142 728 145 738
rect 438 728 441 738
rect 606 728 609 738
rect 806 728 814 731
rect 69 718 70 722
rect 266 718 267 722
rect 388 718 390 722
rect 766 721 769 728
rect 758 718 769 721
rect 680 703 682 707
rect 686 703 689 707
rect 693 703 696 707
rect 738 688 739 692
rect 306 678 313 681
rect 330 678 337 681
rect 86 668 105 671
rect 122 668 124 672
rect 526 668 534 671
rect 786 668 793 671
rect 866 668 873 671
rect 78 658 89 661
rect 174 661 177 668
rect 174 658 185 661
rect 214 658 222 661
rect 230 658 238 661
rect 378 658 385 661
rect 582 658 590 661
rect 746 658 761 661
rect 810 658 817 661
rect 950 658 966 661
rect 86 652 89 658
rect 498 648 502 652
rect 690 648 697 651
rect 762 638 763 642
rect 418 618 419 622
rect 581 618 582 622
rect 670 618 686 621
rect 272 603 274 607
rect 278 603 281 607
rect 285 603 288 607
rect 253 588 254 592
rect 877 588 878 592
rect 646 568 657 571
rect 654 562 657 568
rect 230 558 241 561
rect 30 551 34 554
rect 14 548 34 551
rect 206 551 210 554
rect 190 548 210 551
rect 254 548 273 551
rect 382 548 401 551
rect 406 548 414 551
rect 446 551 449 561
rect 430 548 449 551
rect 522 548 529 551
rect 598 548 610 551
rect 630 548 649 551
rect 678 548 694 551
rect 834 548 841 551
rect 134 541 137 548
rect 126 538 137 541
rect 270 541 273 548
rect 598 542 601 548
rect 606 546 610 548
rect 270 538 297 541
rect 326 538 337 541
rect 342 538 361 541
rect 542 538 553 541
rect 574 538 582 541
rect 758 541 761 548
rect 758 538 769 541
rect 890 538 897 541
rect 334 532 337 538
rect 302 528 318 531
rect 680 503 682 507
rect 686 503 689 507
rect 693 503 696 507
rect 290 488 305 491
rect 378 488 379 492
rect 14 468 25 471
rect 150 468 169 471
rect 322 468 337 471
rect 830 471 833 481
rect 830 468 838 471
rect 846 468 854 471
rect 902 468 910 471
rect 950 462 954 464
rect 10 458 17 461
rect 662 458 678 461
rect 906 458 929 461
rect 222 448 241 451
rect 582 448 590 451
rect 638 448 641 458
rect 238 442 241 448
rect 210 418 211 422
rect 272 403 274 407
rect 278 403 281 407
rect 285 403 288 407
rect 386 388 387 392
rect 458 388 459 392
rect 770 388 771 392
rect 853 388 854 392
rect 38 342 41 351
rect 174 348 185 351
rect 254 348 294 351
rect 318 351 321 361
rect 398 358 409 361
rect 302 348 321 351
rect 182 342 185 348
rect 146 338 161 341
rect 230 338 238 341
rect 274 338 289 341
rect 438 341 441 351
rect 450 348 457 351
rect 570 348 577 351
rect 678 351 681 361
rect 678 348 713 351
rect 734 351 737 361
rect 798 358 809 361
rect 926 358 937 361
rect 942 358 950 361
rect 722 348 737 351
rect 854 348 862 351
rect 438 338 449 341
rect 642 338 657 341
rect 126 328 129 338
rect 438 332 441 338
rect 325 318 326 322
rect 741 318 742 322
rect 680 303 682 307
rect 686 303 689 307
rect 693 303 696 307
rect 678 278 705 281
rect 110 268 118 271
rect 158 268 166 271
rect 390 271 393 278
rect 390 268 409 271
rect 626 268 633 271
rect 782 268 790 271
rect 806 271 809 281
rect 894 278 902 282
rect 934 278 945 281
rect 894 272 897 278
rect 806 268 822 271
rect 842 268 849 271
rect 22 258 41 261
rect 78 258 97 261
rect 450 258 473 261
rect 514 258 521 261
rect 646 258 665 261
rect 786 258 793 261
rect 810 258 817 261
rect 78 256 82 258
rect 318 248 329 251
rect 374 248 385 251
rect 838 248 849 251
rect 326 242 329 248
rect 290 238 297 241
rect 229 228 230 232
rect 925 218 926 222
rect 272 203 274 207
rect 278 203 281 207
rect 285 203 288 207
rect 82 168 83 172
rect 150 166 154 168
rect 302 168 329 171
rect 302 166 306 168
rect 74 148 81 151
rect 98 148 105 151
rect 134 151 137 158
rect 214 152 217 161
rect 262 158 270 161
rect 134 148 145 151
rect 154 148 169 151
rect 346 148 353 151
rect 718 148 726 151
rect 742 148 753 151
rect 790 148 798 151
rect 66 138 73 141
rect 174 138 182 141
rect 302 141 305 148
rect 926 142 929 151
rect 294 138 305 141
rect 518 138 526 141
rect 558 138 566 141
rect 762 138 777 141
rect 866 138 873 141
rect 206 128 217 131
rect 390 131 393 138
rect 382 128 393 131
rect 454 128 468 131
rect 570 128 577 131
rect 718 128 729 131
rect 734 128 742 131
rect 854 128 865 131
rect 680 103 682 107
rect 686 103 689 107
rect 693 103 696 107
rect 36 88 38 92
rect 173 88 174 92
rect 429 88 430 92
rect 650 88 651 92
rect 746 78 761 81
rect 54 68 62 71
rect 142 68 158 71
rect 174 68 190 71
rect 302 68 321 71
rect 126 61 129 68
rect 366 62 369 71
rect 430 68 438 71
rect 474 68 481 71
rect 662 68 705 71
rect 118 58 129 61
rect 222 58 249 61
rect 302 58 310 61
rect 342 58 361 61
rect 438 58 449 61
rect 710 61 713 71
rect 734 62 737 71
rect 818 68 825 71
rect 958 68 974 71
rect 710 58 726 61
rect 886 58 897 61
rect 342 52 345 58
rect 118 48 129 51
rect 370 48 377 51
rect 272 3 274 7
rect 278 3 281 7
rect 285 3 288 7
<< m2contact >>
rect 274 803 278 807
rect 281 803 285 807
rect 894 788 898 792
rect 918 788 922 792
rect 950 788 954 792
rect 710 778 714 782
rect 6 768 10 772
rect 102 768 106 772
rect 134 768 138 772
rect 382 768 386 772
rect 398 768 402 772
rect 718 768 722 772
rect 758 768 762 772
rect 110 758 114 762
rect 166 758 170 762
rect 270 758 274 762
rect 654 758 658 762
rect 702 758 706 762
rect 118 748 122 752
rect 126 748 130 752
rect 190 748 194 752
rect 238 748 242 752
rect 254 748 258 752
rect 326 748 330 752
rect 358 748 362 752
rect 374 748 378 752
rect 422 748 426 752
rect 446 748 450 752
rect 502 748 506 752
rect 510 748 514 752
rect 614 748 618 752
rect 646 748 650 752
rect 670 748 674 752
rect 710 748 714 752
rect 742 748 746 752
rect 766 748 770 752
rect 782 748 786 752
rect 838 748 842 752
rect 902 748 906 752
rect 926 748 930 752
rect 966 748 970 752
rect 78 738 82 742
rect 86 738 90 742
rect 150 738 154 742
rect 254 738 258 742
rect 358 738 362 742
rect 438 738 442 742
rect 478 738 482 742
rect 534 738 538 742
rect 550 738 554 742
rect 590 738 594 742
rect 678 738 682 742
rect 790 738 794 742
rect 38 728 42 732
rect 46 728 50 732
rect 110 728 114 732
rect 174 728 178 732
rect 302 728 306 732
rect 342 728 346 732
rect 398 728 402 732
rect 446 728 450 732
rect 486 728 490 732
rect 494 728 498 732
rect 526 728 530 732
rect 622 728 626 732
rect 742 728 746 732
rect 766 728 770 732
rect 814 728 818 732
rect 822 728 826 732
rect 70 718 74 722
rect 102 718 106 722
rect 166 718 170 722
rect 214 718 218 722
rect 262 718 266 722
rect 310 718 314 722
rect 350 718 354 722
rect 390 718 394 722
rect 454 718 458 722
rect 470 718 474 722
rect 598 718 602 722
rect 942 718 946 722
rect 682 703 686 707
rect 689 703 693 707
rect 46 688 50 692
rect 734 688 738 692
rect 814 688 818 692
rect 902 688 906 692
rect 926 688 930 692
rect 54 678 58 682
rect 110 678 114 682
rect 198 678 202 682
rect 238 678 242 682
rect 246 678 250 682
rect 286 678 290 682
rect 302 678 306 682
rect 326 678 330 682
rect 358 678 362 682
rect 398 678 402 682
rect 406 678 410 682
rect 534 678 538 682
rect 622 678 626 682
rect 638 678 642 682
rect 782 678 786 682
rect 806 678 810 682
rect 862 678 866 682
rect 894 678 898 682
rect 934 678 938 682
rect 46 668 50 672
rect 118 668 122 672
rect 166 668 170 672
rect 174 668 178 672
rect 190 668 194 672
rect 430 668 434 672
rect 454 668 458 672
rect 470 668 474 672
rect 510 668 514 672
rect 518 668 522 672
rect 534 668 538 672
rect 550 668 554 672
rect 590 668 594 672
rect 598 668 602 672
rect 630 668 634 672
rect 662 668 666 672
rect 726 668 730 672
rect 750 668 754 672
rect 782 668 786 672
rect 862 668 866 672
rect 878 668 882 672
rect 910 668 914 672
rect 958 668 962 672
rect 38 658 42 662
rect 94 658 98 662
rect 134 658 138 662
rect 222 658 226 662
rect 238 658 242 662
rect 262 658 266 662
rect 302 658 306 662
rect 326 658 330 662
rect 350 658 354 662
rect 374 658 378 662
rect 422 658 426 662
rect 446 658 450 662
rect 462 658 466 662
rect 478 658 482 662
rect 502 658 506 662
rect 558 658 562 662
rect 590 658 594 662
rect 606 658 610 662
rect 622 658 626 662
rect 654 658 658 662
rect 710 658 714 662
rect 742 658 746 662
rect 798 658 802 662
rect 806 658 810 662
rect 822 658 826 662
rect 846 658 850 662
rect 886 658 890 662
rect 918 658 922 662
rect 966 658 970 662
rect 70 648 74 652
rect 86 648 90 652
rect 142 648 146 652
rect 150 648 154 652
rect 174 648 178 652
rect 294 648 298 652
rect 486 648 490 652
rect 502 648 506 652
rect 566 648 570 652
rect 686 648 690 652
rect 742 648 746 652
rect 774 648 778 652
rect 854 648 858 652
rect 942 648 946 652
rect 126 638 130 642
rect 222 638 226 642
rect 382 638 386 642
rect 654 638 658 642
rect 710 638 714 642
rect 758 638 762 642
rect 838 638 842 642
rect 158 628 162 632
rect 438 628 442 632
rect 702 628 706 632
rect 846 628 850 632
rect 214 618 218 622
rect 262 618 266 622
rect 326 618 330 622
rect 350 618 354 622
rect 374 618 378 622
rect 414 618 418 622
rect 534 618 538 622
rect 582 618 586 622
rect 686 618 690 622
rect 950 618 954 622
rect 274 603 278 607
rect 281 603 285 607
rect 54 588 58 592
rect 254 588 258 592
rect 486 588 490 592
rect 734 588 738 592
rect 878 588 882 592
rect 910 588 914 592
rect 942 588 946 592
rect 342 578 346 582
rect 46 568 50 572
rect 222 568 226 572
rect 742 568 746 572
rect 22 558 26 562
rect 142 558 146 562
rect 150 558 154 562
rect 198 558 202 562
rect 310 558 314 562
rect 390 558 394 562
rect 38 548 42 552
rect 70 548 74 552
rect 102 548 106 552
rect 118 548 122 552
rect 134 548 138 552
rect 182 548 186 552
rect 214 548 218 552
rect 286 548 290 552
rect 350 548 354 552
rect 366 548 370 552
rect 414 548 418 552
rect 422 548 426 552
rect 494 558 498 562
rect 518 558 522 562
rect 550 558 554 562
rect 654 558 658 562
rect 726 558 730 562
rect 806 558 810 562
rect 846 558 850 562
rect 862 558 866 562
rect 974 558 978 562
rect 462 548 466 552
rect 518 548 522 552
rect 534 548 538 552
rect 566 548 570 552
rect 582 548 586 552
rect 614 548 618 552
rect 694 548 698 552
rect 702 548 706 552
rect 734 548 738 552
rect 758 548 762 552
rect 774 548 778 552
rect 790 548 794 552
rect 798 548 802 552
rect 814 548 818 552
rect 822 548 826 552
rect 830 548 834 552
rect 878 548 882 552
rect 926 548 930 552
rect 958 548 962 552
rect 6 538 10 542
rect 62 538 66 542
rect 94 538 98 542
rect 158 538 162 542
rect 174 538 178 542
rect 262 538 266 542
rect 374 538 378 542
rect 414 538 418 542
rect 470 538 474 542
rect 510 538 514 542
rect 582 538 586 542
rect 598 538 602 542
rect 638 538 642 542
rect 830 538 834 542
rect 886 538 890 542
rect 918 538 922 542
rect 950 538 954 542
rect 966 538 970 542
rect 334 528 338 532
rect 438 528 442 532
rect 478 528 482 532
rect 502 528 506 532
rect 598 528 602 532
rect 614 528 618 532
rect 654 528 658 532
rect 662 528 666 532
rect 710 528 714 532
rect 718 528 722 532
rect 758 528 762 532
rect 782 528 786 532
rect 854 528 858 532
rect 902 528 906 532
rect 86 518 90 522
rect 102 518 106 522
rect 166 518 170 522
rect 446 518 450 522
rect 590 518 594 522
rect 670 518 674 522
rect 682 503 686 507
rect 689 503 693 507
rect 38 488 42 492
rect 70 488 74 492
rect 102 488 106 492
rect 246 488 250 492
rect 286 488 290 492
rect 374 488 378 492
rect 470 488 474 492
rect 502 488 506 492
rect 558 488 562 492
rect 710 488 714 492
rect 902 488 906 492
rect 974 488 978 492
rect 118 478 122 482
rect 126 478 130 482
rect 134 478 138 482
rect 190 478 194 482
rect 462 478 466 482
rect 550 478 554 482
rect 718 478 722 482
rect 6 468 10 472
rect 46 468 50 472
rect 78 468 82 472
rect 182 468 186 472
rect 198 468 202 472
rect 278 468 282 472
rect 318 468 322 472
rect 350 468 354 472
rect 366 468 370 472
rect 398 468 402 472
rect 414 468 418 472
rect 438 468 442 472
rect 454 468 458 472
rect 486 468 490 472
rect 494 468 498 472
rect 510 468 514 472
rect 526 468 530 472
rect 542 468 546 472
rect 566 468 570 472
rect 614 468 618 472
rect 638 468 642 472
rect 646 468 650 472
rect 702 468 706 472
rect 758 468 762 472
rect 774 468 778 472
rect 814 468 818 472
rect 838 478 842 482
rect 902 478 906 482
rect 838 468 842 472
rect 854 468 858 472
rect 910 468 914 472
rect 6 458 10 462
rect 54 458 58 462
rect 86 458 90 462
rect 110 458 114 462
rect 158 458 162 462
rect 206 458 210 462
rect 238 458 242 462
rect 326 458 330 462
rect 358 458 362 462
rect 390 458 394 462
rect 406 458 410 462
rect 422 458 426 462
rect 446 458 450 462
rect 478 458 482 462
rect 534 458 538 462
rect 574 458 578 462
rect 590 458 594 462
rect 606 458 610 462
rect 622 458 626 462
rect 638 458 642 462
rect 654 458 658 462
rect 678 458 682 462
rect 694 458 698 462
rect 734 458 738 462
rect 782 458 786 462
rect 790 458 794 462
rect 806 458 810 462
rect 830 458 834 462
rect 854 458 858 462
rect 894 458 898 462
rect 902 458 906 462
rect 950 458 954 462
rect 958 458 962 462
rect 38 448 42 452
rect 70 448 74 452
rect 262 448 266 452
rect 270 448 274 452
rect 302 448 306 452
rect 382 448 386 452
rect 430 448 434 452
rect 518 448 522 452
rect 590 448 594 452
rect 670 448 674 452
rect 726 448 730 452
rect 798 448 802 452
rect 166 438 170 442
rect 238 438 242 442
rect 246 438 250 442
rect 598 438 602 442
rect 742 438 746 442
rect 766 438 770 442
rect 942 438 946 442
rect 750 428 754 432
rect 134 418 138 422
rect 206 418 210 422
rect 334 418 338 422
rect 502 418 506 422
rect 274 403 278 407
rect 281 403 285 407
rect 382 388 386 392
rect 438 388 442 392
rect 454 388 458 392
rect 766 388 770 392
rect 854 388 858 392
rect 870 388 874 392
rect 470 368 474 372
rect 526 368 530 372
rect 806 368 810 372
rect 30 358 34 362
rect 118 358 122 362
rect 310 358 314 362
rect 14 348 18 352
rect 54 348 58 352
rect 70 348 74 352
rect 86 348 90 352
rect 102 348 106 352
rect 142 348 146 352
rect 214 348 218 352
rect 246 348 250 352
rect 294 348 298 352
rect 542 358 546 362
rect 342 348 346 352
rect 382 348 386 352
rect 6 338 10 342
rect 38 338 42 342
rect 46 338 50 342
rect 62 338 66 342
rect 78 338 82 342
rect 94 338 98 342
rect 126 338 130 342
rect 142 338 146 342
rect 182 338 186 342
rect 190 338 194 342
rect 222 338 226 342
rect 238 338 242 342
rect 270 338 274 342
rect 334 338 338 342
rect 350 338 354 342
rect 374 338 378 342
rect 446 348 450 352
rect 478 348 482 352
rect 502 348 506 352
rect 534 348 538 352
rect 558 348 562 352
rect 566 348 570 352
rect 622 348 626 352
rect 662 348 666 352
rect 702 358 706 362
rect 718 348 722 352
rect 782 358 786 362
rect 838 358 842 362
rect 910 358 914 362
rect 950 358 954 362
rect 766 348 770 352
rect 814 348 818 352
rect 822 348 826 352
rect 862 348 866 352
rect 894 348 898 352
rect 902 348 906 352
rect 510 338 514 342
rect 526 338 530 342
rect 550 338 554 342
rect 566 338 570 342
rect 630 338 634 342
rect 638 338 642 342
rect 670 338 674 342
rect 726 338 730 342
rect 750 338 754 342
rect 758 338 762 342
rect 830 338 834 342
rect 862 338 866 342
rect 878 338 882 342
rect 886 338 890 342
rect 950 338 954 342
rect 150 328 154 332
rect 206 328 210 332
rect 238 328 242 332
rect 262 328 266 332
rect 366 328 370 332
rect 414 328 418 332
rect 422 328 426 332
rect 438 328 442 332
rect 486 328 490 332
rect 494 328 498 332
rect 582 328 586 332
rect 638 328 642 332
rect 790 328 794 332
rect 918 328 922 332
rect 30 318 34 322
rect 118 318 122 322
rect 134 318 138 322
rect 198 318 202 322
rect 326 318 330 322
rect 358 318 362 322
rect 630 318 634 322
rect 742 318 746 322
rect 682 303 686 307
rect 689 303 693 307
rect 158 288 162 292
rect 334 288 338 292
rect 374 288 378 292
rect 582 288 586 292
rect 614 288 618 292
rect 734 288 738 292
rect 798 288 802 292
rect 158 278 162 282
rect 246 278 250 282
rect 310 278 314 282
rect 390 278 394 282
rect 398 278 402 282
rect 462 278 466 282
rect 510 278 514 282
rect 590 278 594 282
rect 622 278 626 282
rect 46 268 50 272
rect 86 268 90 272
rect 118 268 122 272
rect 166 268 170 272
rect 190 268 194 272
rect 206 268 210 272
rect 238 268 242 272
rect 254 268 258 272
rect 350 268 354 272
rect 422 268 426 272
rect 478 268 482 272
rect 494 268 498 272
rect 534 268 538 272
rect 550 268 554 272
rect 574 268 578 272
rect 606 268 610 272
rect 622 268 626 272
rect 726 268 730 272
rect 750 268 754 272
rect 766 268 770 272
rect 790 268 794 272
rect 838 278 842 282
rect 822 268 826 272
rect 838 268 842 272
rect 870 268 874 272
rect 886 268 890 272
rect 894 268 898 272
rect 910 268 914 272
rect 966 268 970 272
rect 62 258 66 262
rect 102 258 106 262
rect 150 258 154 262
rect 198 258 202 262
rect 230 258 234 262
rect 294 258 298 262
rect 334 258 338 262
rect 358 258 362 262
rect 414 258 418 262
rect 430 258 434 262
rect 438 258 442 262
rect 446 258 450 262
rect 502 258 506 262
rect 510 258 514 262
rect 526 258 530 262
rect 542 258 546 262
rect 558 258 562 262
rect 566 258 570 262
rect 598 258 602 262
rect 638 258 642 262
rect 718 258 722 262
rect 774 258 778 262
rect 782 258 786 262
rect 806 258 810 262
rect 862 258 866 262
rect 918 258 922 262
rect 958 258 962 262
rect 30 248 34 252
rect 86 248 90 252
rect 182 248 186 252
rect 214 248 218 252
rect 270 248 274 252
rect 446 248 450 252
rect 654 248 658 252
rect 702 248 706 252
rect 734 248 738 252
rect 758 248 762 252
rect 894 248 898 252
rect 942 248 946 252
rect 6 238 10 242
rect 62 238 66 242
rect 286 238 290 242
rect 326 238 330 242
rect 334 238 338 242
rect 878 238 882 242
rect 230 228 234 232
rect 494 228 498 232
rect 70 218 74 222
rect 662 218 666 222
rect 926 218 930 222
rect 274 203 278 207
rect 281 203 285 207
rect 334 188 338 192
rect 750 188 754 192
rect 902 188 906 192
rect 614 178 618 182
rect 78 168 82 172
rect 94 168 98 172
rect 110 168 114 172
rect 150 168 154 172
rect 470 168 474 172
rect 910 168 914 172
rect 126 158 130 162
rect 134 158 138 162
rect 158 158 162 162
rect 38 148 42 152
rect 70 148 74 152
rect 94 148 98 152
rect 118 148 122 152
rect 270 158 274 162
rect 302 158 306 162
rect 310 158 314 162
rect 366 158 370 162
rect 486 158 490 162
rect 502 158 506 162
rect 558 158 562 162
rect 654 158 658 162
rect 662 158 666 162
rect 798 158 802 162
rect 854 158 858 162
rect 894 158 898 162
rect 150 148 154 152
rect 182 148 186 152
rect 214 148 218 152
rect 230 148 234 152
rect 302 148 306 152
rect 318 148 322 152
rect 342 148 346 152
rect 390 148 394 152
rect 422 148 426 152
rect 430 148 434 152
rect 446 148 450 152
rect 478 148 482 152
rect 494 148 498 152
rect 526 148 530 152
rect 542 148 546 152
rect 590 148 594 152
rect 638 148 642 152
rect 678 148 682 152
rect 726 148 730 152
rect 766 148 770 152
rect 798 148 802 152
rect 814 148 818 152
rect 838 148 842 152
rect 886 148 890 152
rect 902 148 906 152
rect 30 138 34 142
rect 46 138 50 142
rect 62 138 66 142
rect 134 138 138 142
rect 182 138 186 142
rect 190 138 194 142
rect 238 138 242 142
rect 246 138 250 142
rect 286 138 290 142
rect 950 148 954 152
rect 342 138 346 142
rect 390 138 394 142
rect 414 138 418 142
rect 438 138 442 142
rect 502 138 506 142
rect 526 138 530 142
rect 534 138 538 142
rect 566 138 570 142
rect 582 138 586 142
rect 630 138 634 142
rect 686 138 690 142
rect 710 138 714 142
rect 758 138 762 142
rect 822 138 826 142
rect 830 138 834 142
rect 862 138 866 142
rect 878 138 882 142
rect 926 138 930 142
rect 942 138 946 142
rect 54 128 58 132
rect 198 128 202 132
rect 374 128 378 132
rect 398 128 402 132
rect 566 128 570 132
rect 654 128 658 132
rect 742 128 746 132
rect 790 128 794 132
rect 926 128 930 132
rect 262 118 266 122
rect 366 118 370 122
rect 406 118 410 122
rect 662 118 666 122
rect 798 118 802 122
rect 682 103 686 107
rect 689 103 693 107
rect 38 88 42 92
rect 86 88 90 92
rect 126 88 130 92
rect 174 88 178 92
rect 190 88 194 92
rect 430 88 434 92
rect 446 88 450 92
rect 502 88 506 92
rect 606 88 610 92
rect 646 88 650 92
rect 750 88 754 92
rect 766 88 770 92
rect 838 88 842 92
rect 854 88 858 92
rect 934 88 938 92
rect 94 78 98 82
rect 230 78 234 82
rect 310 78 314 82
rect 398 78 402 82
rect 862 78 866 82
rect 902 78 906 82
rect 6 68 10 72
rect 62 68 66 72
rect 102 68 106 72
rect 126 68 130 72
rect 158 68 162 72
rect 190 68 194 72
rect 206 68 210 72
rect 238 68 242 72
rect 254 68 258 72
rect 270 68 274 72
rect 334 68 338 72
rect 70 58 74 62
rect 390 68 394 72
rect 414 68 418 72
rect 438 68 442 72
rect 462 66 466 70
rect 470 68 474 72
rect 526 68 530 72
rect 582 68 586 72
rect 630 68 634 72
rect 646 68 650 72
rect 150 58 154 62
rect 182 58 186 62
rect 214 58 218 62
rect 262 58 266 62
rect 294 58 298 62
rect 310 58 314 62
rect 326 58 330 62
rect 366 58 370 62
rect 406 58 410 62
rect 534 58 538 62
rect 558 58 562 62
rect 638 58 642 62
rect 670 58 674 62
rect 718 68 722 72
rect 774 68 778 72
rect 790 68 794 72
rect 814 68 818 72
rect 910 68 914 72
rect 974 68 978 72
rect 726 58 730 62
rect 734 58 738 62
rect 782 58 786 62
rect 806 58 810 62
rect 846 58 850 62
rect 190 48 194 52
rect 342 48 346 52
rect 350 48 354 52
rect 366 48 370 52
rect 694 48 698 52
rect 750 48 754 52
rect 798 48 802 52
rect 838 48 842 52
rect 550 18 554 22
rect 574 18 578 22
rect 870 18 874 22
rect 274 3 278 7
rect 281 3 285 7
<< metal2 >>
rect 102 828 106 832
rect 326 828 330 832
rect 350 831 354 832
rect 350 828 361 831
rect 102 772 105 828
rect 272 803 274 807
rect 278 803 281 807
rect 285 803 288 807
rect 6 762 9 768
rect 134 762 137 768
rect 170 758 174 761
rect 266 758 270 761
rect 90 738 94 741
rect 46 732 49 738
rect 78 732 81 738
rect 110 732 113 758
rect 118 752 121 758
rect 166 752 169 758
rect 190 752 193 758
rect 254 752 257 758
rect 326 752 329 828
rect 358 752 361 828
rect 470 828 474 832
rect 494 828 498 832
rect 886 831 890 832
rect 910 831 914 832
rect 958 831 962 832
rect 886 828 897 831
rect 910 828 921 831
rect 398 772 401 778
rect 386 768 390 771
rect 374 752 377 768
rect 426 748 430 751
rect 126 732 129 748
rect 238 742 241 748
rect 154 738 158 741
rect 250 738 254 741
rect 174 732 177 738
rect 302 732 305 748
rect 326 742 329 748
rect 342 732 345 748
rect 358 732 361 738
rect 374 732 377 748
rect 398 732 401 738
rect 114 728 118 731
rect 38 691 41 728
rect 162 718 166 721
rect 70 692 73 718
rect 38 688 46 691
rect 50 688 54 691
rect 102 682 105 718
rect 214 712 217 718
rect 194 678 198 681
rect 46 672 49 678
rect 38 602 41 658
rect 54 592 57 678
rect 86 652 89 658
rect 70 642 73 648
rect 6 542 9 568
rect 10 538 14 541
rect 6 472 9 478
rect 6 342 9 458
rect 22 432 25 558
rect 38 492 41 548
rect 46 532 49 568
rect 74 548 78 551
rect 94 542 97 658
rect 66 538 70 541
rect 70 492 73 528
rect 86 512 89 518
rect 94 492 97 538
rect 102 532 105 548
rect 110 532 113 678
rect 122 668 126 671
rect 186 668 190 671
rect 130 658 134 661
rect 142 652 145 658
rect 150 642 153 648
rect 126 632 129 638
rect 158 632 161 638
rect 118 552 121 578
rect 142 562 145 568
rect 150 552 153 558
rect 134 542 137 548
rect 154 538 158 541
rect 166 532 169 668
rect 174 662 177 668
rect 222 662 225 698
rect 238 692 241 728
rect 238 682 241 688
rect 246 682 249 688
rect 262 672 265 718
rect 286 682 289 728
rect 302 682 305 718
rect 310 702 313 718
rect 350 682 353 718
rect 358 682 361 718
rect 326 672 329 678
rect 262 662 265 668
rect 302 662 305 668
rect 326 662 329 668
rect 350 662 353 678
rect 374 662 377 698
rect 390 692 393 718
rect 406 682 409 748
rect 438 732 441 738
rect 446 732 449 748
rect 470 732 473 828
rect 494 752 497 828
rect 894 792 897 828
rect 918 792 921 828
rect 950 828 962 831
rect 950 792 953 828
rect 710 762 713 778
rect 722 768 726 771
rect 762 768 766 771
rect 646 752 649 758
rect 498 748 502 751
rect 478 742 481 748
rect 482 728 486 731
rect 498 728 502 731
rect 510 722 513 748
rect 590 742 593 748
rect 538 738 542 741
rect 530 728 534 731
rect 394 678 398 681
rect 422 662 425 678
rect 454 672 457 718
rect 470 681 473 718
rect 470 678 478 681
rect 242 658 246 661
rect 174 622 177 648
rect 222 642 225 648
rect 214 622 217 628
rect 214 612 217 618
rect 254 592 257 598
rect 262 591 265 618
rect 272 603 274 607
rect 278 603 281 607
rect 285 603 288 607
rect 262 588 273 591
rect 222 562 225 568
rect 202 558 209 561
rect 174 532 177 538
rect 102 512 105 518
rect 106 488 110 491
rect 118 482 121 528
rect 134 492 137 528
rect 158 492 161 518
rect 166 512 169 518
rect 134 482 137 488
rect 114 478 118 481
rect 46 472 49 478
rect 126 472 129 478
rect 82 468 86 471
rect 158 462 161 488
rect 182 482 185 548
rect 206 522 209 558
rect 214 542 217 548
rect 190 472 193 478
rect 198 472 201 478
rect 46 451 49 458
rect 42 448 49 451
rect 54 452 57 458
rect 86 452 89 458
rect 110 452 113 458
rect 182 452 185 468
rect 206 462 209 518
rect 246 492 249 538
rect 262 502 265 538
rect 270 492 273 588
rect 286 492 289 548
rect 238 462 241 488
rect 274 468 278 471
rect 274 448 278 451
rect 14 352 17 408
rect 34 358 38 361
rect 38 342 41 348
rect 46 342 49 448
rect 70 442 73 448
rect 54 352 57 358
rect 70 352 73 408
rect 86 352 89 388
rect 82 348 86 351
rect 94 342 97 358
rect 6 332 9 338
rect 30 261 33 318
rect 62 312 65 338
rect 50 268 54 271
rect 62 262 65 298
rect 30 258 41 261
rect 6 242 9 248
rect 30 242 33 248
rect 30 142 33 238
rect 38 152 41 258
rect 58 238 62 241
rect 70 222 73 228
rect 78 211 81 338
rect 94 332 97 338
rect 102 332 105 348
rect 110 332 113 448
rect 170 438 174 441
rect 182 422 185 448
rect 238 442 241 448
rect 250 438 254 441
rect 262 422 265 448
rect 294 432 297 648
rect 378 638 382 641
rect 430 632 433 668
rect 442 658 446 661
rect 462 652 465 658
rect 442 628 446 631
rect 330 618 334 621
rect 378 618 385 621
rect 350 612 353 618
rect 350 592 353 608
rect 342 572 345 578
rect 314 558 318 561
rect 310 512 313 558
rect 350 552 353 558
rect 354 548 361 551
rect 334 532 337 548
rect 338 528 342 531
rect 350 472 353 528
rect 358 482 361 548
rect 366 542 369 548
rect 374 542 377 568
rect 382 512 385 618
rect 398 562 401 618
rect 390 522 393 558
rect 374 492 377 498
rect 318 452 321 468
rect 358 462 361 478
rect 302 442 305 448
rect 326 442 329 458
rect 294 422 297 428
rect 118 362 121 368
rect 134 352 137 418
rect 206 382 209 418
rect 272 403 274 407
rect 278 403 281 407
rect 285 403 288 407
rect 146 358 153 361
rect 142 352 145 358
rect 126 332 129 338
rect 142 332 145 338
rect 150 332 153 358
rect 90 268 94 271
rect 102 262 105 278
rect 118 272 121 318
rect 134 262 137 318
rect 158 292 161 298
rect 154 278 158 281
rect 150 262 153 268
rect 86 242 89 248
rect 70 208 81 211
rect 70 152 73 208
rect 94 192 97 258
rect 94 172 97 188
rect 78 162 81 168
rect 50 138 54 141
rect 50 128 54 131
rect 38 92 41 108
rect 6 72 9 88
rect 62 72 65 138
rect 70 92 73 148
rect 94 132 97 148
rect 102 132 105 258
rect 158 252 161 278
rect 166 272 169 358
rect 182 342 185 348
rect 190 342 193 368
rect 246 352 249 388
rect 334 382 337 418
rect 366 372 369 468
rect 382 452 385 508
rect 390 462 393 478
rect 398 472 401 558
rect 414 552 417 618
rect 438 572 441 628
rect 470 562 473 668
rect 478 662 481 678
rect 502 662 505 708
rect 534 682 537 688
rect 550 672 553 738
rect 594 718 598 721
rect 530 668 534 671
rect 482 648 486 651
rect 502 642 505 648
rect 510 602 513 668
rect 518 612 521 668
rect 486 582 489 588
rect 490 558 494 561
rect 466 548 470 551
rect 422 542 425 548
rect 510 542 513 598
rect 534 562 537 618
rect 522 558 526 561
rect 522 548 526 551
rect 414 512 417 538
rect 410 468 414 471
rect 398 462 401 468
rect 422 462 425 488
rect 438 472 441 528
rect 446 502 449 518
rect 454 472 457 518
rect 470 492 473 538
rect 498 528 502 531
rect 478 492 481 528
rect 502 492 505 518
rect 446 462 449 468
rect 382 392 385 428
rect 306 358 310 361
rect 210 348 214 351
rect 290 348 294 351
rect 338 348 342 351
rect 234 338 238 341
rect 190 332 193 338
rect 222 332 225 338
rect 234 328 238 331
rect 194 318 198 321
rect 206 312 209 328
rect 246 282 249 348
rect 350 342 353 358
rect 342 338 350 341
rect 254 328 262 331
rect 254 272 257 328
rect 270 322 273 338
rect 186 268 190 271
rect 210 268 214 271
rect 242 268 246 271
rect 150 172 153 238
rect 110 162 113 168
rect 126 162 129 168
rect 134 152 137 158
rect 150 152 153 158
rect 158 152 161 158
rect 122 148 126 151
rect 86 92 89 98
rect 126 92 129 128
rect 134 102 137 138
rect 166 122 169 268
rect 194 258 198 261
rect 226 258 230 261
rect 174 248 182 251
rect 210 248 214 251
rect 70 62 73 88
rect 94 72 97 78
rect 102 72 105 88
rect 158 72 161 98
rect 174 92 177 248
rect 234 228 238 231
rect 182 152 185 158
rect 190 142 193 168
rect 214 152 217 158
rect 230 152 233 168
rect 254 142 257 268
rect 294 262 297 318
rect 310 282 313 288
rect 326 272 329 318
rect 334 292 337 338
rect 318 258 326 261
rect 330 258 334 261
rect 274 248 278 251
rect 282 238 286 241
rect 272 203 274 207
rect 278 203 281 207
rect 285 203 288 207
rect 270 162 273 178
rect 302 162 305 168
rect 250 138 254 141
rect 182 82 185 138
rect 198 122 201 128
rect 190 92 193 118
rect 214 72 217 118
rect 230 82 233 138
rect 238 112 241 138
rect 238 72 241 88
rect 254 72 257 128
rect 270 122 273 158
rect 302 142 305 148
rect 262 102 265 118
rect 286 112 289 138
rect 310 112 313 158
rect 318 152 321 258
rect 326 242 329 248
rect 334 232 337 238
rect 342 212 345 338
rect 366 322 369 328
rect 358 282 361 318
rect 374 311 377 338
rect 366 308 377 311
rect 382 312 385 348
rect 398 322 401 458
rect 406 452 409 458
rect 422 352 425 458
rect 430 452 433 458
rect 454 392 457 408
rect 462 392 465 478
rect 486 472 489 478
rect 510 472 513 508
rect 498 468 502 471
rect 482 458 486 461
rect 518 461 521 508
rect 534 502 537 548
rect 542 491 545 668
rect 534 488 545 491
rect 550 662 553 668
rect 558 662 561 708
rect 590 672 593 678
rect 550 562 553 658
rect 558 648 566 651
rect 550 492 553 558
rect 558 492 561 648
rect 582 552 585 618
rect 590 592 593 658
rect 598 632 601 668
rect 606 662 609 728
rect 614 642 617 748
rect 654 742 657 758
rect 622 722 625 728
rect 670 722 673 748
rect 678 732 681 738
rect 680 703 682 707
rect 686 703 689 707
rect 693 703 696 707
rect 626 678 630 681
rect 634 678 638 681
rect 658 668 662 671
rect 622 662 625 668
rect 630 662 633 668
rect 646 658 654 661
rect 646 652 649 658
rect 682 648 686 651
rect 654 642 657 648
rect 598 612 601 628
rect 614 552 617 608
rect 686 592 689 618
rect 654 562 657 568
rect 694 552 697 678
rect 702 662 705 758
rect 714 748 718 751
rect 738 748 742 751
rect 762 748 766 751
rect 906 748 910 751
rect 782 742 785 748
rect 838 742 841 748
rect 742 722 745 728
rect 766 722 769 728
rect 734 692 737 698
rect 742 672 745 718
rect 782 712 785 738
rect 790 732 793 738
rect 806 682 809 708
rect 814 692 817 728
rect 822 722 825 728
rect 814 682 817 688
rect 786 678 790 681
rect 750 672 753 678
rect 778 668 782 671
rect 710 651 713 658
rect 726 652 729 668
rect 742 662 745 668
rect 846 662 849 708
rect 862 682 865 698
rect 902 692 905 738
rect 926 692 929 748
rect 894 682 897 688
rect 942 682 945 718
rect 878 672 881 678
rect 866 668 870 671
rect 906 668 910 671
rect 878 658 886 661
rect 710 648 721 651
rect 734 648 742 651
rect 718 642 721 648
rect 734 642 737 648
rect 758 642 761 648
rect 702 632 705 638
rect 710 612 713 638
rect 734 592 737 638
rect 746 568 750 571
rect 726 562 729 568
rect 702 552 705 558
rect 570 548 574 551
rect 598 542 601 548
rect 586 538 590 541
rect 638 532 641 538
rect 654 532 657 538
rect 602 528 606 531
rect 618 528 622 531
rect 662 522 665 528
rect 694 521 697 548
rect 702 542 705 548
rect 718 532 721 548
rect 734 542 737 548
rect 758 542 761 548
rect 706 528 710 531
rect 766 531 769 658
rect 774 652 777 658
rect 798 602 801 658
rect 762 528 769 531
rect 774 552 777 588
rect 806 562 809 658
rect 814 552 817 608
rect 822 592 825 658
rect 834 638 838 641
rect 846 632 849 648
rect 854 622 857 648
rect 822 552 825 558
rect 830 552 833 598
rect 878 592 881 658
rect 918 652 921 658
rect 934 622 937 678
rect 942 652 945 668
rect 958 652 961 668
rect 966 662 969 748
rect 910 592 913 598
rect 942 592 945 598
rect 862 562 865 568
rect 842 558 846 561
rect 786 548 790 551
rect 694 518 713 521
rect 590 502 593 518
rect 526 472 529 478
rect 510 458 521 461
rect 534 462 537 488
rect 546 478 550 481
rect 442 388 446 391
rect 470 372 473 398
rect 478 352 481 368
rect 502 362 505 418
rect 498 348 502 351
rect 438 332 441 338
rect 446 332 449 348
rect 510 342 513 458
rect 522 448 526 451
rect 526 372 529 378
rect 534 362 537 458
rect 542 442 545 468
rect 566 422 569 468
rect 590 462 593 488
rect 614 472 617 488
rect 638 472 641 478
rect 578 458 585 461
rect 602 458 606 461
rect 566 382 569 418
rect 542 362 545 368
rect 558 352 561 358
rect 582 352 585 458
rect 590 402 593 448
rect 602 438 606 441
rect 590 372 593 398
rect 614 392 617 468
rect 626 458 630 461
rect 638 452 641 458
rect 646 442 649 468
rect 654 462 657 468
rect 670 452 673 518
rect 680 503 682 507
rect 686 503 689 507
rect 693 503 696 507
rect 710 492 713 518
rect 718 472 721 478
rect 682 458 686 461
rect 694 452 697 458
rect 702 412 705 468
rect 734 462 737 478
rect 750 472 753 528
rect 774 482 777 548
rect 782 532 785 538
rect 798 522 801 548
rect 822 538 830 541
rect 754 468 758 471
rect 770 468 774 471
rect 810 468 814 471
rect 726 452 729 458
rect 742 442 745 458
rect 762 438 766 441
rect 750 422 753 428
rect 766 392 769 408
rect 638 388 646 391
rect 538 348 542 351
rect 570 348 574 351
rect 522 338 526 341
rect 546 338 550 341
rect 410 328 414 331
rect 426 328 430 331
rect 366 302 369 308
rect 374 292 377 298
rect 350 262 353 268
rect 358 252 361 258
rect 330 188 334 191
rect 274 68 278 71
rect 126 62 129 68
rect 146 58 150 61
rect 182 52 185 58
rect 190 52 193 68
rect 206 52 209 68
rect 214 62 217 68
rect 294 62 297 78
rect 310 72 313 78
rect 326 62 329 98
rect 334 72 337 168
rect 342 152 345 208
rect 366 162 369 198
rect 382 172 385 308
rect 390 282 393 318
rect 422 302 425 328
rect 478 322 481 338
rect 486 322 489 328
rect 494 322 497 328
rect 390 242 393 258
rect 362 158 366 161
rect 390 152 393 238
rect 398 172 401 278
rect 462 272 465 278
rect 478 272 481 318
rect 510 282 513 308
rect 526 302 529 338
rect 550 272 553 318
rect 566 302 569 338
rect 574 302 577 348
rect 582 332 585 348
rect 622 342 625 348
rect 638 342 641 388
rect 698 358 702 361
rect 774 361 777 468
rect 790 462 793 468
rect 822 462 825 538
rect 850 528 854 531
rect 834 478 838 481
rect 850 468 854 471
rect 826 458 830 461
rect 782 402 785 458
rect 798 452 801 458
rect 806 372 809 458
rect 838 442 841 468
rect 850 458 854 461
rect 774 358 782 361
rect 630 332 633 338
rect 642 328 646 331
rect 426 268 430 271
rect 418 258 422 261
rect 450 258 454 261
rect 430 252 433 258
rect 438 222 441 258
rect 430 152 433 188
rect 446 152 449 248
rect 422 142 425 148
rect 342 102 345 138
rect 390 132 393 138
rect 414 132 417 138
rect 366 122 369 128
rect 374 92 377 128
rect 398 122 401 128
rect 410 118 414 121
rect 266 58 270 61
rect 306 58 310 61
rect 342 52 345 58
rect 350 52 353 78
rect 390 72 393 78
rect 398 72 401 78
rect 366 62 369 68
rect 406 62 409 108
rect 430 92 433 138
rect 438 122 441 138
rect 450 88 454 91
rect 462 82 465 268
rect 494 242 497 268
rect 526 262 529 268
rect 514 258 518 261
rect 502 252 505 258
rect 534 252 537 268
rect 542 252 545 258
rect 498 228 502 231
rect 470 142 473 168
rect 478 152 481 228
rect 486 162 489 168
rect 494 152 497 178
rect 502 162 505 168
rect 510 151 513 248
rect 542 152 545 208
rect 502 148 513 151
rect 522 148 526 151
rect 502 142 505 148
rect 502 92 505 98
rect 526 92 529 138
rect 534 132 537 138
rect 442 68 446 71
rect 462 70 465 78
rect 526 72 529 78
rect 414 52 417 68
rect 470 62 473 68
rect 534 62 537 98
rect 550 82 553 268
rect 558 262 561 298
rect 614 292 617 318
rect 586 288 590 291
rect 622 282 625 288
rect 594 278 598 281
rect 602 268 606 271
rect 618 268 622 271
rect 566 262 569 268
rect 566 161 569 258
rect 574 192 577 268
rect 594 258 598 261
rect 562 158 569 161
rect 582 142 585 218
rect 614 182 617 188
rect 630 162 633 318
rect 638 262 641 268
rect 654 262 657 358
rect 714 348 718 351
rect 662 342 665 348
rect 718 342 721 348
rect 670 332 673 338
rect 726 332 729 338
rect 750 332 753 338
rect 680 303 682 307
rect 686 303 689 307
rect 693 303 696 307
rect 742 302 745 318
rect 758 312 761 338
rect 766 332 769 348
rect 786 328 790 331
rect 738 288 742 291
rect 730 268 737 271
rect 714 258 718 261
rect 646 248 654 251
rect 698 248 702 251
rect 590 152 593 158
rect 630 142 633 148
rect 638 142 641 148
rect 570 138 574 141
rect 626 138 630 141
rect 566 122 569 128
rect 566 61 569 118
rect 582 102 585 138
rect 638 92 641 138
rect 646 92 649 248
rect 654 162 657 198
rect 662 162 665 218
rect 726 152 729 268
rect 734 252 737 268
rect 750 242 753 268
rect 758 252 761 298
rect 766 272 769 328
rect 798 292 801 368
rect 814 352 817 398
rect 838 362 841 438
rect 854 392 857 418
rect 862 412 865 558
rect 874 548 878 551
rect 886 532 889 538
rect 902 532 905 538
rect 902 492 905 508
rect 902 462 905 478
rect 910 472 913 558
rect 918 542 921 578
rect 950 562 953 618
rect 954 548 958 551
rect 918 522 921 538
rect 926 512 929 548
rect 950 482 953 538
rect 894 452 897 458
rect 870 392 873 448
rect 902 432 905 458
rect 942 442 945 448
rect 858 348 862 351
rect 822 282 825 348
rect 830 332 833 338
rect 838 282 841 348
rect 878 342 881 348
rect 886 342 889 368
rect 894 352 897 378
rect 950 372 953 458
rect 958 382 961 458
rect 914 358 918 361
rect 946 358 950 361
rect 902 352 905 358
rect 950 342 953 348
rect 862 322 865 338
rect 826 268 830 271
rect 750 192 753 228
rect 678 132 681 148
rect 758 142 761 148
rect 766 142 769 148
rect 714 138 718 141
rect 686 132 689 138
rect 738 128 742 131
rect 654 122 657 128
rect 666 118 670 121
rect 562 58 569 61
rect 610 88 614 91
rect 582 72 585 88
rect 642 68 646 71
rect 370 48 374 51
rect 190 42 193 48
rect 350 22 353 48
rect 366 42 369 48
rect 272 3 274 7
rect 278 3 281 7
rect 285 3 288 7
rect 334 -18 337 18
rect 470 -18 473 58
rect 334 -22 338 -18
rect 470 -22 474 -18
rect 542 -19 546 -18
rect 550 -19 553 18
rect 542 -22 553 -19
rect 566 -19 570 -18
rect 574 -19 577 18
rect 582 12 585 68
rect 630 52 633 68
rect 670 62 673 108
rect 680 103 682 107
rect 686 103 689 107
rect 693 103 696 107
rect 750 92 753 118
rect 766 92 769 128
rect 774 122 777 258
rect 782 142 785 258
rect 790 242 793 268
rect 794 158 798 161
rect 794 148 798 151
rect 806 132 809 258
rect 838 162 841 268
rect 862 262 865 278
rect 870 272 873 328
rect 886 272 889 338
rect 922 328 926 331
rect 894 272 897 278
rect 890 248 894 251
rect 850 158 854 161
rect 818 148 822 151
rect 830 142 833 148
rect 838 142 841 148
rect 870 142 873 248
rect 878 232 881 238
rect 902 192 905 328
rect 910 272 913 278
rect 918 262 921 318
rect 966 282 969 538
rect 974 492 977 558
rect 910 172 913 178
rect 926 162 929 218
rect 882 148 886 151
rect 874 138 878 141
rect 822 132 825 138
rect 642 58 646 61
rect 694 52 697 78
rect 722 68 726 71
rect 718 52 721 68
rect 734 62 737 68
rect 774 62 777 68
rect 782 62 785 78
rect 790 72 793 128
rect 802 118 806 121
rect 854 92 857 128
rect 842 88 846 91
rect 862 82 865 138
rect 894 132 897 158
rect 906 148 910 151
rect 902 82 905 148
rect 926 142 929 148
rect 926 122 929 128
rect 934 92 937 268
rect 942 252 945 258
rect 942 142 945 158
rect 950 152 953 278
rect 962 268 966 271
rect 962 258 966 261
rect 910 72 913 78
rect 974 72 977 258
rect 786 58 790 61
rect 726 52 729 58
rect 566 -22 577 -19
rect 630 -18 633 48
rect 750 12 753 48
rect 774 42 777 58
rect 806 52 809 58
rect 794 48 798 51
rect 814 12 817 68
rect 846 62 849 68
rect 838 42 841 48
rect 734 -18 737 8
rect 630 -22 634 -18
rect 734 -22 738 -18
rect 870 -19 873 18
rect 934 -18 937 8
rect 878 -19 882 -18
rect 870 -22 882 -19
rect 934 -22 938 -18
<< m3contact >>
rect 274 803 278 807
rect 281 803 285 807
rect 6 758 10 762
rect 118 758 122 762
rect 134 758 138 762
rect 174 758 178 762
rect 190 758 194 762
rect 254 758 258 762
rect 262 758 266 762
rect 46 738 50 742
rect 94 738 98 742
rect 398 778 402 782
rect 374 768 378 772
rect 390 768 394 772
rect 166 748 170 752
rect 302 748 306 752
rect 342 748 346 752
rect 358 748 362 752
rect 406 748 410 752
rect 430 748 434 752
rect 158 738 162 742
rect 174 738 178 742
rect 238 738 242 742
rect 246 738 250 742
rect 326 738 330 742
rect 398 738 402 742
rect 78 728 82 732
rect 118 728 122 732
rect 126 728 130 732
rect 238 728 242 732
rect 286 728 290 732
rect 358 728 362 732
rect 374 728 378 732
rect 158 718 162 722
rect 54 688 58 692
rect 70 688 74 692
rect 214 708 218 712
rect 222 698 226 702
rect 46 678 50 682
rect 102 678 106 682
rect 190 678 194 682
rect 38 598 42 602
rect 86 658 90 662
rect 70 638 74 642
rect 6 568 10 572
rect 14 538 18 542
rect 6 478 10 482
rect 78 548 82 552
rect 70 538 74 542
rect 46 528 50 532
rect 70 528 74 532
rect 86 508 90 512
rect 126 668 130 672
rect 182 668 186 672
rect 126 658 130 662
rect 142 658 146 662
rect 150 638 154 642
rect 158 638 162 642
rect 126 628 130 632
rect 118 578 122 582
rect 142 568 146 572
rect 150 548 154 552
rect 134 538 138 542
rect 150 538 154 542
rect 238 688 242 692
rect 246 688 250 692
rect 302 718 306 722
rect 358 718 362 722
rect 310 698 314 702
rect 374 698 378 702
rect 350 678 354 682
rect 262 668 266 672
rect 302 668 306 672
rect 326 668 330 672
rect 390 688 394 692
rect 726 768 730 772
rect 766 768 770 772
rect 646 758 650 762
rect 710 758 714 762
rect 478 748 482 752
rect 494 748 498 752
rect 590 748 594 752
rect 438 728 442 732
rect 470 728 474 732
rect 478 728 482 732
rect 502 728 506 732
rect 542 738 546 742
rect 534 728 538 732
rect 454 718 458 722
rect 510 718 514 722
rect 390 678 394 682
rect 422 678 426 682
rect 502 708 506 712
rect 478 678 482 682
rect 174 658 178 662
rect 246 658 250 662
rect 222 648 226 652
rect 214 628 218 632
rect 174 618 178 622
rect 262 618 266 622
rect 214 608 218 612
rect 254 598 258 602
rect 274 603 278 607
rect 281 603 285 607
rect 198 558 202 562
rect 222 558 226 562
rect 102 528 106 532
rect 110 528 114 532
rect 118 528 122 532
rect 134 528 138 532
rect 166 528 170 532
rect 174 528 178 532
rect 102 508 106 512
rect 94 488 98 492
rect 110 488 114 492
rect 158 518 162 522
rect 166 508 170 512
rect 134 488 138 492
rect 158 488 162 492
rect 46 478 50 482
rect 110 478 114 482
rect 86 468 90 472
rect 126 468 130 472
rect 214 538 218 542
rect 246 538 250 542
rect 206 518 210 522
rect 182 478 186 482
rect 198 478 202 482
rect 190 468 194 472
rect 46 458 50 462
rect 262 498 266 502
rect 238 488 242 492
rect 270 488 274 492
rect 270 468 274 472
rect 54 448 58 452
rect 86 448 90 452
rect 110 448 114 452
rect 182 448 186 452
rect 238 448 242 452
rect 278 448 282 452
rect 22 428 26 432
rect 14 408 18 412
rect 38 358 42 362
rect 38 348 42 352
rect 70 438 74 442
rect 70 408 74 412
rect 54 358 58 362
rect 86 388 90 392
rect 94 358 98 362
rect 78 348 82 352
rect 78 338 82 342
rect 6 328 10 332
rect 62 308 66 312
rect 62 298 66 302
rect 54 268 58 272
rect 6 248 10 252
rect 30 238 34 242
rect 54 238 58 242
rect 70 228 74 232
rect 174 438 178 442
rect 254 438 258 442
rect 374 638 378 642
rect 438 658 442 662
rect 462 648 466 652
rect 430 628 434 632
rect 446 628 450 632
rect 334 618 338 622
rect 350 608 354 612
rect 350 588 354 592
rect 342 568 346 572
rect 374 568 378 572
rect 318 558 322 562
rect 350 558 354 562
rect 334 548 338 552
rect 342 528 346 532
rect 350 528 354 532
rect 310 508 314 512
rect 366 538 370 542
rect 398 618 402 622
rect 398 558 402 562
rect 390 518 394 522
rect 382 508 386 512
rect 374 498 378 502
rect 358 478 362 482
rect 318 448 322 452
rect 302 438 306 442
rect 326 438 330 442
rect 294 428 298 432
rect 182 418 186 422
rect 262 418 266 422
rect 294 418 298 422
rect 118 368 122 372
rect 274 403 278 407
rect 281 403 285 407
rect 246 388 250 392
rect 206 378 210 382
rect 190 368 194 372
rect 142 358 146 362
rect 134 348 138 352
rect 166 358 170 362
rect 94 328 98 332
rect 102 328 106 332
rect 110 328 114 332
rect 126 328 130 332
rect 142 328 146 332
rect 102 278 106 282
rect 94 268 98 272
rect 158 298 162 302
rect 150 278 154 282
rect 150 268 154 272
rect 94 258 98 262
rect 134 258 138 262
rect 86 238 90 242
rect 94 188 98 192
rect 78 158 82 162
rect 54 138 58 142
rect 62 138 66 142
rect 46 128 50 132
rect 38 108 42 112
rect 6 88 10 92
rect 182 348 186 352
rect 334 378 338 382
rect 390 478 394 482
rect 438 568 442 572
rect 534 688 538 692
rect 606 728 610 732
rect 590 718 594 722
rect 558 708 562 712
rect 526 668 530 672
rect 542 668 546 672
rect 478 648 482 652
rect 502 638 506 642
rect 518 608 522 612
rect 510 598 514 602
rect 486 578 490 582
rect 470 558 474 562
rect 486 558 490 562
rect 470 548 474 552
rect 526 558 530 562
rect 534 558 538 562
rect 526 548 530 552
rect 422 538 426 542
rect 414 508 418 512
rect 422 488 426 492
rect 406 468 410 472
rect 454 518 458 522
rect 446 498 450 502
rect 494 528 498 532
rect 502 518 506 522
rect 510 508 514 512
rect 518 508 522 512
rect 478 488 482 492
rect 486 478 490 482
rect 446 468 450 472
rect 398 458 402 462
rect 430 458 434 462
rect 382 428 386 432
rect 366 368 370 372
rect 302 358 306 362
rect 350 358 354 362
rect 206 348 210 352
rect 286 348 290 352
rect 334 348 338 352
rect 230 338 234 342
rect 190 328 194 332
rect 222 328 226 332
rect 230 328 234 332
rect 190 318 194 322
rect 206 308 210 312
rect 270 318 274 322
rect 294 318 298 322
rect 182 268 186 272
rect 214 268 218 272
rect 246 268 250 272
rect 158 248 162 252
rect 150 238 154 242
rect 126 168 130 172
rect 110 158 114 162
rect 150 158 154 162
rect 126 148 130 152
rect 134 148 138 152
rect 158 148 162 152
rect 94 128 98 132
rect 102 128 106 132
rect 126 128 130 132
rect 86 98 90 102
rect 190 258 194 262
rect 222 258 226 262
rect 206 248 210 252
rect 166 118 170 122
rect 134 98 138 102
rect 158 98 162 102
rect 70 88 74 92
rect 102 88 106 92
rect 62 68 66 72
rect 238 228 242 232
rect 190 168 194 172
rect 230 168 234 172
rect 182 158 186 162
rect 214 158 218 162
rect 310 288 314 292
rect 326 268 330 272
rect 326 258 330 262
rect 278 248 282 252
rect 278 238 282 242
rect 274 203 278 207
rect 281 203 285 207
rect 270 178 274 182
rect 302 168 306 172
rect 230 138 234 142
rect 254 138 258 142
rect 190 118 194 122
rect 198 118 202 122
rect 214 118 218 122
rect 182 78 186 82
rect 254 128 258 132
rect 238 108 242 112
rect 238 88 242 92
rect 302 138 306 142
rect 270 118 274 122
rect 326 248 330 252
rect 334 228 338 232
rect 366 318 370 322
rect 406 448 410 452
rect 454 408 458 412
rect 502 468 506 472
rect 486 458 490 462
rect 534 498 538 502
rect 590 678 594 682
rect 550 658 554 662
rect 654 738 658 742
rect 678 728 682 732
rect 622 718 626 722
rect 670 718 674 722
rect 682 703 686 707
rect 689 703 693 707
rect 630 678 634 682
rect 694 678 698 682
rect 622 668 626 672
rect 654 668 658 672
rect 630 658 634 662
rect 646 648 650 652
rect 654 648 658 652
rect 678 648 682 652
rect 614 638 618 642
rect 598 628 602 632
rect 598 608 602 612
rect 614 608 618 612
rect 590 588 594 592
rect 686 588 690 592
rect 654 568 658 572
rect 718 748 722 752
rect 734 748 738 752
rect 758 748 762 752
rect 910 748 914 752
rect 966 748 970 752
rect 782 738 786 742
rect 838 738 842 742
rect 902 738 906 742
rect 742 718 746 722
rect 766 718 770 722
rect 734 698 738 702
rect 790 728 794 732
rect 782 708 786 712
rect 806 708 810 712
rect 822 718 826 722
rect 846 708 850 712
rect 750 678 754 682
rect 790 678 794 682
rect 814 678 818 682
rect 742 668 746 672
rect 774 668 778 672
rect 702 658 706 662
rect 862 698 866 702
rect 894 688 898 692
rect 878 678 882 682
rect 942 678 946 682
rect 870 668 874 672
rect 902 668 906 672
rect 766 658 770 662
rect 774 658 778 662
rect 726 648 730 652
rect 758 648 762 652
rect 702 638 706 642
rect 718 638 722 642
rect 734 638 738 642
rect 710 608 714 612
rect 726 568 730 572
rect 750 568 754 572
rect 702 558 706 562
rect 574 548 578 552
rect 598 548 602 552
rect 718 548 722 552
rect 590 538 594 542
rect 654 538 658 542
rect 606 528 610 532
rect 622 528 626 532
rect 638 528 642 532
rect 662 518 666 522
rect 702 538 706 542
rect 734 538 738 542
rect 758 538 762 542
rect 702 528 706 532
rect 750 528 754 532
rect 798 598 802 602
rect 774 588 778 592
rect 814 608 818 612
rect 846 648 850 652
rect 830 638 834 642
rect 854 618 858 622
rect 830 598 834 602
rect 822 588 826 592
rect 822 558 826 562
rect 918 648 922 652
rect 942 668 946 672
rect 958 648 962 652
rect 934 618 938 622
rect 910 598 914 602
rect 942 598 946 602
rect 918 578 922 582
rect 862 568 866 572
rect 838 558 842 562
rect 910 558 914 562
rect 782 548 786 552
rect 830 548 834 552
rect 590 498 594 502
rect 550 488 554 492
rect 590 488 594 492
rect 614 488 618 492
rect 526 478 530 482
rect 542 478 546 482
rect 470 398 474 402
rect 446 388 450 392
rect 462 388 466 392
rect 478 368 482 372
rect 502 358 506 362
rect 422 348 426 352
rect 494 348 498 352
rect 438 338 442 342
rect 526 448 530 452
rect 526 378 530 382
rect 542 438 546 442
rect 638 478 642 482
rect 654 468 658 472
rect 598 458 602 462
rect 566 418 570 422
rect 566 378 570 382
rect 542 368 546 372
rect 534 358 538 362
rect 558 358 562 362
rect 606 438 610 442
rect 590 398 594 402
rect 630 458 634 462
rect 638 448 642 452
rect 682 503 686 507
rect 689 503 693 507
rect 734 478 738 482
rect 718 468 722 472
rect 686 458 690 462
rect 694 448 698 452
rect 646 438 650 442
rect 782 538 786 542
rect 798 518 802 522
rect 774 478 778 482
rect 750 468 754 472
rect 766 468 770 472
rect 790 468 794 472
rect 806 468 810 472
rect 726 458 730 462
rect 742 458 746 462
rect 758 438 762 442
rect 750 418 754 422
rect 702 408 706 412
rect 766 408 770 412
rect 614 388 618 392
rect 646 388 650 392
rect 590 368 594 372
rect 542 348 546 352
rect 574 348 578 352
rect 582 348 586 352
rect 478 338 482 342
rect 518 338 522 342
rect 542 338 546 342
rect 406 328 410 332
rect 430 328 434 332
rect 446 328 450 332
rect 390 318 394 322
rect 398 318 402 322
rect 382 308 386 312
rect 366 298 370 302
rect 374 298 378 302
rect 358 278 362 282
rect 350 258 354 262
rect 358 248 362 252
rect 342 208 346 212
rect 326 188 330 192
rect 334 168 338 172
rect 286 108 290 112
rect 310 108 314 112
rect 262 98 266 102
rect 326 98 330 102
rect 294 78 298 82
rect 94 68 98 72
rect 102 68 106 72
rect 214 68 218 72
rect 278 68 282 72
rect 126 58 130 62
rect 142 58 146 62
rect 310 68 314 72
rect 366 198 370 202
rect 478 318 482 322
rect 486 318 490 322
rect 494 318 498 322
rect 422 298 426 302
rect 390 258 394 262
rect 390 238 394 242
rect 382 168 386 172
rect 358 158 362 162
rect 510 308 514 312
rect 550 318 554 322
rect 526 298 530 302
rect 654 358 658 362
rect 694 358 698 362
rect 846 528 850 532
rect 830 478 834 482
rect 846 468 850 472
rect 798 458 802 462
rect 822 458 826 462
rect 782 398 786 402
rect 846 458 850 462
rect 838 438 842 442
rect 814 398 818 402
rect 798 368 802 372
rect 622 338 626 342
rect 630 328 634 332
rect 646 328 650 332
rect 614 318 618 322
rect 558 298 562 302
rect 566 298 570 302
rect 574 298 578 302
rect 430 268 434 272
rect 462 268 466 272
rect 526 268 530 272
rect 422 258 426 262
rect 454 258 458 262
rect 430 248 434 252
rect 438 218 442 222
rect 430 188 434 192
rect 398 168 402 172
rect 422 138 426 142
rect 430 138 434 142
rect 366 128 370 132
rect 390 128 394 132
rect 414 128 418 132
rect 342 98 346 102
rect 398 118 402 122
rect 414 118 418 122
rect 406 108 410 112
rect 374 88 378 92
rect 350 78 354 82
rect 390 78 394 82
rect 270 58 274 62
rect 302 58 306 62
rect 342 58 346 62
rect 366 68 370 72
rect 398 68 402 72
rect 438 118 442 122
rect 454 88 458 92
rect 518 258 522 262
rect 502 248 506 252
rect 510 248 514 252
rect 534 248 538 252
rect 542 248 546 252
rect 494 238 498 242
rect 478 228 482 232
rect 502 228 506 232
rect 494 178 498 182
rect 486 168 490 172
rect 502 168 506 172
rect 542 208 546 212
rect 518 148 522 152
rect 470 138 474 142
rect 502 98 506 102
rect 534 128 538 132
rect 534 98 538 102
rect 526 88 530 92
rect 462 78 466 82
rect 526 78 530 82
rect 446 68 450 72
rect 590 288 594 292
rect 622 288 626 292
rect 598 278 602 282
rect 566 268 570 272
rect 598 268 602 272
rect 614 268 618 272
rect 590 258 594 262
rect 582 218 586 222
rect 574 188 578 192
rect 614 188 618 192
rect 638 268 642 272
rect 710 348 714 352
rect 662 338 666 342
rect 718 338 722 342
rect 670 328 674 332
rect 726 328 730 332
rect 750 328 754 332
rect 682 303 686 307
rect 689 303 693 307
rect 766 328 770 332
rect 782 328 786 332
rect 758 308 762 312
rect 742 298 746 302
rect 758 298 762 302
rect 742 288 746 292
rect 654 258 658 262
rect 710 258 714 262
rect 694 248 698 252
rect 590 158 594 162
rect 630 158 634 162
rect 630 148 634 152
rect 574 138 578 142
rect 622 138 626 142
rect 638 138 642 142
rect 566 118 570 122
rect 550 78 554 82
rect 470 58 474 62
rect 582 98 586 102
rect 654 198 658 202
rect 854 418 858 422
rect 870 548 874 552
rect 902 538 906 542
rect 886 528 890 532
rect 902 508 906 512
rect 950 558 954 562
rect 950 548 954 552
rect 918 518 922 522
rect 926 508 930 512
rect 950 478 954 482
rect 870 448 874 452
rect 894 448 898 452
rect 862 408 866 412
rect 942 448 946 452
rect 902 428 906 432
rect 894 378 898 382
rect 886 368 890 372
rect 838 348 842 352
rect 854 348 858 352
rect 878 348 882 352
rect 830 328 834 332
rect 958 378 962 382
rect 950 368 954 372
rect 902 358 906 362
rect 918 358 922 362
rect 942 358 946 362
rect 950 348 954 352
rect 870 328 874 332
rect 862 318 866 322
rect 822 278 826 282
rect 862 278 866 282
rect 830 268 834 272
rect 750 238 754 242
rect 750 228 754 232
rect 758 148 762 152
rect 718 138 722 142
rect 766 138 770 142
rect 678 128 682 132
rect 686 128 690 132
rect 734 128 738 132
rect 766 128 770 132
rect 654 118 658 122
rect 670 118 674 122
rect 750 118 754 122
rect 670 108 674 112
rect 582 88 586 92
rect 614 88 618 92
rect 638 88 642 92
rect 638 68 642 72
rect 182 48 186 52
rect 206 48 210 52
rect 374 48 378 52
rect 414 48 418 52
rect 190 38 194 42
rect 366 38 370 42
rect 334 18 338 22
rect 350 18 354 22
rect 274 3 278 7
rect 281 3 285 7
rect 682 103 686 107
rect 689 103 693 107
rect 790 238 794 242
rect 790 158 794 162
rect 790 148 794 152
rect 782 138 786 142
rect 902 328 906 332
rect 926 328 930 332
rect 894 278 898 282
rect 886 268 890 272
rect 870 248 874 252
rect 886 248 890 252
rect 838 158 842 162
rect 846 158 850 162
rect 822 148 826 152
rect 830 148 834 152
rect 878 228 882 232
rect 918 318 922 322
rect 910 278 914 282
rect 950 278 954 282
rect 966 278 970 282
rect 934 268 938 272
rect 910 178 914 182
rect 926 158 930 162
rect 878 148 882 152
rect 838 138 842 142
rect 870 138 874 142
rect 806 128 810 132
rect 822 128 826 132
rect 854 128 858 132
rect 774 118 778 122
rect 766 88 770 92
rect 694 78 698 82
rect 782 78 786 82
rect 646 58 650 62
rect 726 68 730 72
rect 734 68 738 72
rect 806 118 810 122
rect 846 88 850 92
rect 910 148 914 152
rect 926 148 930 152
rect 894 128 898 132
rect 926 118 930 122
rect 942 258 946 262
rect 942 158 946 162
rect 958 268 962 272
rect 966 258 970 262
rect 974 258 978 262
rect 910 78 914 82
rect 846 68 850 72
rect 774 58 778 62
rect 790 58 794 62
rect 630 48 634 52
rect 718 48 722 52
rect 726 48 730 52
rect 582 8 586 12
rect 790 48 794 52
rect 806 48 810 52
rect 774 38 778 42
rect 838 38 842 42
rect 734 8 738 12
rect 750 8 754 12
rect 814 8 818 12
rect 934 8 938 12
<< metal3 >>
rect 272 803 274 807
rect 278 803 281 807
rect 286 803 288 807
rect 134 768 374 771
rect 398 771 401 778
rect 394 768 401 771
rect 730 768 758 771
rect 762 768 766 771
rect 134 762 137 768
rect -26 761 -22 762
rect -26 758 6 761
rect 178 758 190 761
rect 258 758 262 761
rect 650 758 710 761
rect 118 751 121 758
rect 118 748 166 751
rect 306 748 342 751
rect 346 748 358 751
rect 362 748 406 751
rect 434 748 478 751
rect 482 748 494 751
rect 498 748 590 751
rect 722 748 734 751
rect 738 748 758 751
rect 914 748 966 751
rect -26 741 -22 742
rect -26 738 46 741
rect 50 738 94 741
rect 98 738 158 741
rect 162 738 174 741
rect 242 738 246 741
rect 250 738 326 741
rect 330 738 398 741
rect 546 738 654 741
rect 658 738 782 741
rect 842 738 902 741
rect 790 732 793 738
rect 82 728 118 731
rect 122 728 126 731
rect 242 728 286 731
rect 362 728 374 731
rect 442 728 470 731
rect 474 728 478 731
rect 506 728 534 731
rect 538 728 606 731
rect 682 728 702 731
rect 622 722 625 728
rect 822 722 825 728
rect 162 718 302 721
rect 306 718 358 721
rect 458 718 510 721
rect 594 718 614 721
rect 674 718 742 721
rect 770 718 817 721
rect 42 708 214 711
rect 218 708 470 711
rect 474 708 502 711
rect 670 711 673 718
rect 562 708 673 711
rect 786 708 806 711
rect 814 711 817 718
rect 814 708 846 711
rect 680 703 682 707
rect 686 703 689 707
rect 694 703 696 707
rect 226 698 310 701
rect 314 698 374 701
rect 738 698 862 701
rect 50 688 54 691
rect 74 688 238 691
rect 394 688 534 691
rect 590 688 894 691
rect 106 678 190 681
rect 246 681 249 688
rect 590 682 593 688
rect 194 678 249 681
rect 354 678 390 681
rect 394 678 422 681
rect 482 678 590 681
rect 622 678 630 681
rect 698 678 702 681
rect 706 678 750 681
rect 786 678 790 681
rect 818 678 878 681
rect 938 678 942 681
rect 46 671 49 678
rect 46 668 126 671
rect 186 668 190 671
rect 266 668 302 671
rect 306 668 326 671
rect 530 668 542 671
rect 546 668 622 671
rect 658 668 662 671
rect 746 668 774 671
rect 874 668 902 671
rect 906 668 942 671
rect 90 658 126 661
rect 146 658 174 661
rect 250 658 438 661
rect 554 658 630 661
rect 634 658 702 661
rect 706 658 766 661
rect 770 658 774 661
rect 154 648 222 651
rect 466 648 478 651
rect 502 648 646 651
rect 658 648 678 651
rect 682 648 726 651
rect 850 648 918 651
rect 922 648 958 651
rect 70 642 73 648
rect 150 642 153 648
rect 502 642 505 648
rect 226 638 374 641
rect 618 638 702 641
rect 722 638 734 641
rect 758 641 761 648
rect 758 638 830 641
rect 158 631 161 638
rect 130 628 161 631
rect 218 628 430 631
rect 450 628 598 631
rect 178 618 262 621
rect 338 618 398 621
rect 514 618 790 621
rect 794 618 846 621
rect 850 618 854 621
rect 906 618 934 621
rect 82 608 214 611
rect 354 608 478 611
rect 482 608 518 611
rect 602 608 614 611
rect 714 608 814 611
rect 272 603 274 607
rect 278 603 281 607
rect 286 603 288 607
rect 42 598 254 601
rect 514 598 798 601
rect 802 598 830 601
rect 834 598 910 601
rect 1006 601 1010 602
rect 946 598 1010 601
rect 74 588 350 591
rect 486 588 590 591
rect 594 588 614 591
rect 690 588 774 591
rect 778 588 822 591
rect 486 582 489 588
rect 122 578 345 581
rect 1006 581 1010 582
rect 922 578 1010 581
rect 342 572 345 578
rect -26 571 -22 572
rect -26 568 6 571
rect 378 568 438 571
rect 658 568 726 571
rect 754 568 862 571
rect 142 561 145 568
rect 222 562 225 568
rect 142 558 198 561
rect 322 558 350 561
rect 402 558 470 561
rect 474 558 486 561
rect 530 558 534 561
rect 706 558 822 561
rect 826 558 838 561
rect 914 558 950 561
rect 1006 561 1010 562
rect 978 558 1010 561
rect -26 551 -22 552
rect -26 548 78 551
rect 82 548 150 551
rect 154 548 334 551
rect 366 548 425 551
rect 474 548 526 551
rect 578 548 598 551
rect 602 548 718 551
rect 722 548 782 551
rect 834 548 870 551
rect 954 548 958 551
rect 366 542 369 548
rect 422 542 425 548
rect 18 538 70 541
rect 74 538 134 541
rect 138 538 150 541
rect 218 538 246 541
rect 594 538 654 541
rect 658 538 702 541
rect 738 538 758 541
rect 786 538 902 541
rect 906 538 974 541
rect 782 532 785 538
rect 50 528 70 531
rect 106 528 110 531
rect 114 528 118 531
rect 138 528 166 531
rect 170 528 174 531
rect 346 528 350 531
rect 498 528 518 531
rect 610 528 622 531
rect 642 528 646 531
rect 706 528 750 531
rect 850 528 886 531
rect 86 518 158 521
rect 210 518 390 521
rect 394 518 454 521
rect 506 518 622 521
rect 626 518 662 521
rect 670 518 798 521
rect 802 518 918 521
rect 86 512 89 518
rect 106 508 110 511
rect 170 508 310 511
rect 386 508 414 511
rect 418 508 510 511
rect 670 511 673 518
rect 522 508 673 511
rect 906 508 926 511
rect 680 503 682 507
rect 686 503 689 507
rect 694 503 696 507
rect 266 498 374 501
rect 450 498 454 501
rect 538 498 542 501
rect 594 498 670 501
rect 98 488 110 491
rect 114 488 134 491
rect 162 488 238 491
rect 274 488 422 491
rect 426 488 478 491
rect 554 488 590 491
rect 618 488 889 491
rect 886 482 889 488
rect 114 478 182 481
rect 186 478 198 481
rect 362 478 390 481
rect 442 478 486 481
rect 530 478 542 481
rect 674 478 734 481
rect 778 478 830 481
rect 834 478 838 481
rect 890 478 950 481
rect -26 471 -22 472
rect 6 471 9 478
rect 46 471 49 478
rect -26 468 86 471
rect 90 468 126 471
rect 130 468 190 471
rect 194 468 270 471
rect 274 468 406 471
rect 450 468 502 471
rect 506 468 630 471
rect 638 471 641 478
rect 638 468 654 471
rect 722 468 750 471
rect 754 468 766 471
rect 810 468 814 471
rect 826 468 846 471
rect 50 458 398 461
rect 490 458 598 461
rect 602 458 609 461
rect 626 458 630 461
rect 690 458 726 461
rect 790 461 793 468
rect 746 458 793 461
rect 802 458 814 461
rect 826 458 846 461
rect -26 451 -22 452
rect -26 448 54 451
rect 58 448 86 451
rect 90 448 110 451
rect 114 448 182 451
rect 242 448 278 451
rect 282 448 318 451
rect 430 451 433 458
rect 894 452 897 458
rect 410 448 433 451
rect 522 448 526 451
rect 538 448 638 451
rect 642 448 694 451
rect 698 448 870 451
rect 1006 451 1010 452
rect 946 448 1010 451
rect 74 438 78 441
rect 178 438 254 441
rect 258 438 302 441
rect 306 438 326 441
rect 546 438 606 441
rect 610 438 646 441
rect 650 438 758 441
rect 762 438 838 441
rect 382 432 385 438
rect 26 428 294 431
rect 750 428 902 431
rect 750 422 753 428
rect 186 418 262 421
rect 298 418 566 421
rect 762 418 854 421
rect 70 412 73 418
rect 18 408 38 411
rect 458 408 702 411
rect 770 408 862 411
rect 272 403 274 407
rect 278 403 281 407
rect 286 403 288 407
rect 474 398 590 401
rect 786 398 814 401
rect 90 388 246 391
rect 450 388 462 391
rect 466 388 614 391
rect 642 388 646 391
rect 210 378 230 381
rect 242 378 334 381
rect 538 378 566 381
rect 898 378 950 381
rect 954 378 958 381
rect 106 368 118 371
rect 122 368 190 371
rect 194 368 366 371
rect 474 368 478 371
rect 526 371 529 378
rect 526 368 542 371
rect 594 368 798 371
rect 890 368 950 371
rect 42 358 54 361
rect 98 358 142 361
rect 170 358 302 361
rect 306 358 350 361
rect 434 358 502 361
rect 538 358 558 361
rect 562 358 654 361
rect 674 358 694 361
rect 922 358 942 361
rect 42 348 78 351
rect 138 348 142 351
rect 186 348 206 351
rect 290 348 334 351
rect 426 348 494 351
rect 498 348 502 351
rect 546 348 574 351
rect 586 348 710 351
rect 834 348 838 351
rect 858 348 878 351
rect 902 351 905 358
rect 882 348 905 351
rect 82 338 190 341
rect 234 338 438 341
rect 482 338 518 341
rect 546 338 622 341
rect 666 338 702 341
rect 722 338 910 341
rect 950 341 953 348
rect 1006 341 1010 342
rect 914 338 1010 341
rect 10 328 94 331
rect 106 328 110 331
rect 114 328 126 331
rect 130 328 142 331
rect 194 328 222 331
rect 234 328 246 331
rect 410 328 414 331
rect 434 328 446 331
rect 486 328 630 331
rect 650 328 670 331
rect 730 328 750 331
rect 754 328 758 331
rect 770 328 782 331
rect 826 328 830 331
rect 834 328 870 331
rect 898 328 902 331
rect 922 328 926 331
rect 486 322 489 328
rect 194 318 270 321
rect 274 318 294 321
rect 370 318 390 321
rect 402 318 478 321
rect 498 318 550 321
rect 618 318 862 321
rect 866 318 918 321
rect 66 308 190 311
rect 194 308 206 311
rect 386 308 510 311
rect 730 308 758 311
rect 680 303 682 307
rect 686 303 689 307
rect 694 303 696 307
rect 50 298 62 301
rect 162 298 366 301
rect 378 298 422 301
rect 530 298 558 301
rect 578 298 622 301
rect 706 298 742 301
rect 746 298 758 301
rect 566 292 569 298
rect 314 288 430 291
rect 582 288 590 291
rect 594 288 598 291
rect 626 288 630 291
rect 634 288 742 291
rect 106 278 150 281
rect 362 278 422 281
rect 450 278 598 281
rect 602 278 822 281
rect 826 278 862 281
rect 866 278 894 281
rect 954 278 966 281
rect 430 272 433 278
rect 58 268 94 271
rect 146 268 150 271
rect 186 268 198 271
rect 218 268 238 271
rect 242 268 246 271
rect 330 268 382 271
rect 466 268 526 271
rect 602 268 606 271
rect 618 268 622 271
rect 834 268 886 271
rect 910 271 913 278
rect 890 268 934 271
rect 938 268 958 271
rect 82 258 94 261
rect 138 258 190 261
rect 194 258 222 261
rect 330 258 350 261
rect 354 258 390 261
rect 426 258 454 261
rect 482 258 505 261
rect 566 261 569 268
rect 522 258 569 261
rect 594 258 598 261
rect 638 261 641 268
rect 618 258 641 261
rect 658 258 710 261
rect 850 258 942 261
rect 954 258 966 261
rect 1006 261 1010 262
rect 978 258 1010 261
rect 502 252 505 258
rect -26 251 -22 252
rect -26 248 6 251
rect 162 248 206 251
rect 282 248 326 251
rect 330 248 358 251
rect 386 248 430 251
rect 514 248 534 251
rect 546 248 694 251
rect 874 248 886 251
rect 890 248 958 251
rect 86 242 89 248
rect 150 242 153 248
rect 34 238 54 241
rect 162 238 278 241
rect 394 238 494 241
rect 498 238 502 241
rect 570 238 750 241
rect 754 238 790 241
rect 794 238 798 241
rect 802 238 881 241
rect 878 232 881 238
rect 230 228 238 231
rect 242 228 334 231
rect 482 228 502 231
rect 754 228 830 231
rect 70 221 73 228
rect 70 218 430 221
rect 442 218 582 221
rect 346 208 542 211
rect 272 203 274 207
rect 278 203 281 207
rect 286 203 288 207
rect 370 198 654 201
rect 658 198 662 201
rect 98 188 318 191
rect 330 188 430 191
rect 434 188 574 191
rect 274 178 494 181
rect 614 181 617 188
rect 614 178 910 181
rect 230 172 233 178
rect 78 168 113 171
rect 78 162 81 168
rect 110 162 113 168
rect 194 168 230 171
rect 234 168 302 171
rect 338 168 382 171
rect 126 161 129 168
rect 398 162 401 168
rect 126 158 150 161
rect 186 158 190 161
rect 218 158 222 161
rect 226 158 358 161
rect 486 161 489 168
rect 502 161 505 168
rect 846 162 849 168
rect 486 158 505 161
rect 634 158 790 161
rect 826 158 838 161
rect 930 158 942 161
rect 590 152 593 158
rect 130 148 134 151
rect 162 148 494 151
rect 498 148 518 151
rect 634 148 758 151
rect 794 148 822 151
rect 834 148 878 151
rect 882 148 886 151
rect 914 148 926 151
rect 50 138 54 141
rect 66 138 230 141
rect 234 138 254 141
rect 306 138 422 141
rect 434 138 470 141
rect 578 138 622 141
rect 642 138 718 141
rect 722 138 766 141
rect 770 138 782 141
rect 786 138 838 141
rect 842 138 870 141
rect 50 128 94 131
rect 106 128 126 131
rect 138 128 201 131
rect 250 128 254 131
rect 394 128 414 131
rect 422 131 425 138
rect 422 128 534 131
rect 654 128 678 131
rect 690 128 734 131
rect 770 128 806 131
rect 826 128 830 131
rect 858 128 894 131
rect 898 128 902 131
rect 198 122 201 128
rect 170 118 190 121
rect 218 118 270 121
rect 366 121 369 128
rect 654 122 657 128
rect 366 118 398 121
rect 406 118 414 121
rect 418 118 438 121
rect 458 118 566 121
rect 662 118 670 121
rect 674 118 742 121
rect 754 118 774 121
rect 798 118 806 121
rect 810 118 926 121
rect 42 108 182 111
rect 186 108 238 111
rect 242 108 286 111
rect 290 108 310 111
rect 322 108 406 111
rect 410 108 670 111
rect 680 103 682 107
rect 686 103 689 107
rect 694 103 696 107
rect 90 98 134 101
rect 162 98 262 101
rect 266 98 326 101
rect 330 98 342 101
rect 538 98 582 101
rect -26 91 -22 92
rect -26 88 6 91
rect 10 88 70 91
rect 74 88 102 91
rect 134 91 137 98
rect 502 92 505 98
rect 134 88 238 91
rect 242 88 374 91
rect 386 88 454 91
rect 530 88 582 91
rect 618 88 638 91
rect 650 88 766 91
rect 850 88 950 91
rect 186 78 294 81
rect 298 78 350 81
rect 354 78 390 81
rect 394 78 462 81
rect 466 78 526 81
rect 554 78 694 81
rect 698 78 782 81
rect 910 72 913 78
rect -26 71 -22 72
rect -26 68 62 71
rect 66 68 94 71
rect 106 68 214 71
rect 274 68 278 71
rect 314 68 366 71
rect 370 68 398 71
rect 442 68 446 71
rect 450 68 638 71
rect 730 68 734 71
rect 746 68 846 71
rect 130 58 142 61
rect 274 58 302 61
rect 398 61 401 68
rect 398 58 470 61
rect 650 58 654 61
rect 726 58 774 61
rect 794 58 809 61
rect 186 48 206 51
rect 342 51 345 58
rect 726 52 729 58
rect 806 52 809 58
rect 210 48 345 51
rect 378 48 414 51
rect 634 48 718 51
rect 794 48 798 51
rect 194 38 366 41
rect 778 38 838 41
rect 338 18 350 21
rect 586 8 734 11
rect 738 8 750 11
rect 754 8 814 11
rect 938 8 942 11
rect 272 3 274 7
rect 278 3 281 7
rect 286 3 288 7
<< m4contact >>
rect 274 803 278 807
rect 282 803 285 807
rect 285 803 286 807
rect 758 768 762 772
rect 790 738 794 742
rect 622 728 626 732
rect 702 728 706 732
rect 822 728 826 732
rect 614 718 618 722
rect 38 708 42 712
rect 470 708 474 712
rect 682 703 686 707
rect 690 703 693 707
rect 693 703 694 707
rect 46 688 50 692
rect 702 678 706 682
rect 782 678 786 682
rect 934 678 938 682
rect 190 668 194 672
rect 662 668 666 672
rect 438 658 442 662
rect 70 648 74 652
rect 150 648 154 652
rect 222 638 226 642
rect 510 618 514 622
rect 790 618 794 622
rect 846 618 850 622
rect 902 618 906 622
rect 78 608 82 612
rect 478 608 482 612
rect 274 603 278 607
rect 282 603 285 607
rect 285 603 286 607
rect 70 588 74 592
rect 614 588 618 592
rect 222 568 226 572
rect 974 558 978 562
rect 958 548 962 552
rect 974 538 978 542
rect 518 528 522 532
rect 646 528 650 532
rect 782 528 786 532
rect 622 518 626 522
rect 110 508 114 512
rect 510 508 514 512
rect 682 503 686 507
rect 690 503 693 507
rect 693 503 694 507
rect 454 498 458 502
rect 542 498 546 502
rect 670 498 674 502
rect 438 478 442 482
rect 670 478 674 482
rect 838 478 842 482
rect 886 478 890 482
rect 630 468 634 472
rect 814 468 818 472
rect 822 468 826 472
rect 622 458 626 462
rect 814 458 818 462
rect 894 458 898 462
rect 518 448 522 452
rect 534 448 538 452
rect 78 438 82 442
rect 382 438 386 442
rect 70 418 74 422
rect 758 418 762 422
rect 38 408 42 412
rect 274 403 278 407
rect 282 403 285 407
rect 285 403 286 407
rect 638 388 642 392
rect 230 378 234 382
rect 238 378 242 382
rect 534 378 538 382
rect 950 378 954 382
rect 102 368 106 372
rect 470 368 474 372
rect 430 358 434 362
rect 670 358 674 362
rect 142 348 146 352
rect 502 348 506 352
rect 830 348 834 352
rect 190 338 194 342
rect 702 338 706 342
rect 910 338 914 342
rect 246 328 250 332
rect 414 328 418 332
rect 758 328 762 332
rect 822 328 826 332
rect 894 328 898 332
rect 918 328 922 332
rect 190 308 194 312
rect 726 308 730 312
rect 682 303 686 307
rect 690 303 693 307
rect 693 303 694 307
rect 46 298 50 302
rect 622 298 626 302
rect 702 298 706 302
rect 430 288 434 292
rect 566 288 570 292
rect 598 288 602 292
rect 630 288 634 292
rect 422 278 426 282
rect 430 278 434 282
rect 446 278 450 282
rect 142 268 146 272
rect 198 268 202 272
rect 238 268 242 272
rect 382 268 386 272
rect 606 268 610 272
rect 622 268 626 272
rect 78 258 82 262
rect 478 258 482 262
rect 598 258 602 262
rect 614 258 618 262
rect 846 258 850 262
rect 950 258 954 262
rect 974 258 978 262
rect 86 248 90 252
rect 150 248 154 252
rect 382 248 386 252
rect 534 248 538 252
rect 958 248 962 252
rect 158 238 162 242
rect 502 238 506 242
rect 566 238 570 242
rect 798 238 802 242
rect 830 228 834 232
rect 430 218 434 222
rect 274 203 278 207
rect 282 203 285 207
rect 285 203 286 207
rect 662 198 666 202
rect 318 188 322 192
rect 230 178 234 182
rect 846 168 850 172
rect 190 158 194 162
rect 222 158 226 162
rect 398 158 402 162
rect 822 158 826 162
rect 494 148 498 152
rect 590 148 594 152
rect 886 148 890 152
rect 46 138 50 142
rect 134 128 138 132
rect 246 128 250 132
rect 830 128 834 132
rect 902 128 906 132
rect 454 118 458 122
rect 742 118 746 122
rect 182 108 186 112
rect 318 108 322 112
rect 670 108 674 112
rect 682 103 686 107
rect 690 103 693 107
rect 693 103 694 107
rect 382 88 386 92
rect 502 88 506 92
rect 646 88 650 92
rect 950 88 954 92
rect 270 68 274 72
rect 398 68 402 72
rect 438 68 442 72
rect 742 68 746 72
rect 910 68 914 72
rect 654 58 658 62
rect 798 48 802 52
rect 942 8 946 12
rect 274 3 278 7
rect 282 3 285 7
rect 285 3 286 7
<< metal4 >>
rect 272 803 274 807
rect 278 803 281 807
rect 286 803 288 807
rect 614 722 617 728
rect 38 412 41 708
rect 46 302 49 688
rect 70 592 73 648
rect 70 422 73 588
rect 78 442 81 608
rect 102 508 110 511
rect 78 262 81 438
rect 102 372 105 508
rect 142 272 145 348
rect 150 252 153 648
rect 190 342 193 668
rect 222 572 225 638
rect 272 603 274 607
rect 278 603 281 607
rect 286 603 288 607
rect 90 248 94 251
rect 158 242 161 248
rect 190 162 193 308
rect 202 268 206 271
rect 222 162 225 568
rect 438 482 441 658
rect 382 442 385 468
rect 272 403 274 407
rect 278 403 281 407
rect 286 403 288 407
rect 230 182 233 378
rect 238 272 241 378
rect 418 328 422 331
rect 182 158 190 161
rect 50 138 54 141
rect 134 132 137 138
rect 182 112 185 158
rect 246 132 249 328
rect 430 292 433 358
rect 430 282 433 288
rect 382 252 385 268
rect 422 262 425 278
rect 272 203 274 207
rect 278 203 281 207
rect 286 203 288 207
rect 318 112 321 188
rect 382 72 385 88
rect 398 72 401 158
rect 430 152 433 218
rect 438 72 441 478
rect 446 282 449 328
rect 454 122 457 498
rect 470 372 473 708
rect 478 262 481 608
rect 510 512 513 618
rect 518 452 521 528
rect 534 498 542 501
rect 534 452 537 498
rect 494 348 502 351
rect 494 152 497 348
rect 534 252 537 378
rect 602 288 606 291
rect 566 242 569 288
rect 602 268 606 271
rect 614 262 617 588
rect 622 522 625 728
rect 680 703 682 707
rect 686 703 689 707
rect 694 703 696 707
rect 702 682 705 728
rect 638 528 646 531
rect 638 471 641 528
rect 634 468 641 471
rect 626 458 633 461
rect 622 272 625 298
rect 630 292 633 458
rect 638 392 641 468
rect 594 258 598 261
rect 502 92 505 238
rect 662 202 665 668
rect 680 503 682 507
rect 686 503 689 507
rect 694 503 696 507
rect 670 482 673 498
rect 758 422 761 768
rect 782 532 785 678
rect 790 622 793 738
rect 818 728 822 731
rect 810 468 814 471
rect 822 461 825 468
rect 818 458 825 461
rect 586 148 590 151
rect 670 112 673 358
rect 838 351 841 478
rect 834 348 841 351
rect 680 303 682 307
rect 686 303 689 307
rect 694 303 696 307
rect 702 302 705 338
rect 754 328 758 331
rect 826 328 833 331
rect 726 292 729 308
rect 680 103 682 107
rect 686 103 689 107
rect 694 103 696 107
rect 274 68 278 71
rect 646 61 649 88
rect 742 72 745 118
rect 646 58 654 61
rect 798 52 801 238
rect 830 232 833 328
rect 846 262 849 618
rect 846 172 849 258
rect 822 131 825 158
rect 886 152 889 478
rect 894 332 897 458
rect 902 132 905 618
rect 822 128 830 131
rect 910 72 913 338
rect 922 328 926 331
rect 934 11 937 678
rect 950 262 953 378
rect 950 92 953 258
rect 958 252 961 548
rect 974 542 977 558
rect 974 262 977 328
rect 934 8 942 11
rect 272 3 274 7
rect 278 3 281 7
rect 286 3 288 7
<< m5contact >>
rect 274 803 278 807
rect 281 803 282 807
rect 282 803 285 807
rect 614 728 618 732
rect 274 603 278 607
rect 281 603 282 607
rect 282 603 285 607
rect 94 248 98 252
rect 158 248 162 252
rect 206 268 210 272
rect 382 468 386 472
rect 274 403 278 407
rect 281 403 282 407
rect 282 403 285 407
rect 422 328 426 332
rect 54 138 58 142
rect 134 138 138 142
rect 422 258 426 262
rect 274 203 278 207
rect 281 203 282 207
rect 282 203 285 207
rect 430 148 434 152
rect 446 328 450 332
rect 606 288 610 292
rect 598 268 602 272
rect 682 703 686 707
rect 689 703 690 707
rect 690 703 693 707
rect 590 258 594 262
rect 682 503 686 507
rect 689 503 690 507
rect 690 503 693 507
rect 814 728 818 732
rect 806 468 810 472
rect 582 148 586 152
rect 682 303 686 307
rect 689 303 690 307
rect 690 303 693 307
rect 750 328 754 332
rect 726 288 730 292
rect 682 103 686 107
rect 689 103 690 107
rect 690 103 693 107
rect 278 68 282 72
rect 382 68 386 72
rect 926 328 930 332
rect 974 328 978 332
rect 274 3 278 7
rect 281 3 282 7
rect 282 3 285 7
<< metal5 >>
rect 278 803 281 807
rect 277 802 282 803
rect 287 802 288 807
rect 618 728 814 731
rect 686 703 689 707
rect 685 702 690 703
rect 695 702 696 707
rect 278 603 281 607
rect 277 602 282 603
rect 287 602 288 607
rect 686 503 689 507
rect 685 502 690 503
rect 695 502 696 507
rect 386 468 806 471
rect 278 403 281 407
rect 277 402 282 403
rect 287 402 288 407
rect 426 328 446 331
rect 754 328 926 331
rect 930 328 974 331
rect 686 303 689 307
rect 685 302 690 303
rect 695 302 696 307
rect 610 288 726 291
rect 210 268 598 271
rect 426 258 590 261
rect 98 248 158 251
rect 278 203 281 207
rect 277 202 282 203
rect 287 202 288 207
rect 434 148 582 151
rect 58 138 134 141
rect 686 103 689 107
rect 685 102 690 103
rect 695 102 696 107
rect 282 68 382 71
rect 278 3 281 7
rect 277 2 282 3
rect 287 2 288 7
<< m6contact >>
rect 272 803 274 807
rect 274 803 277 807
rect 282 803 285 807
rect 285 803 287 807
rect 272 802 277 803
rect 282 802 287 803
rect 680 703 682 707
rect 682 703 685 707
rect 690 703 693 707
rect 693 703 695 707
rect 680 702 685 703
rect 690 702 695 703
rect 272 603 274 607
rect 274 603 277 607
rect 282 603 285 607
rect 285 603 287 607
rect 272 602 277 603
rect 282 602 287 603
rect 680 503 682 507
rect 682 503 685 507
rect 690 503 693 507
rect 693 503 695 507
rect 680 502 685 503
rect 690 502 695 503
rect 272 403 274 407
rect 274 403 277 407
rect 282 403 285 407
rect 285 403 287 407
rect 272 402 277 403
rect 282 402 287 403
rect 680 303 682 307
rect 682 303 685 307
rect 690 303 693 307
rect 693 303 695 307
rect 680 302 685 303
rect 690 302 695 303
rect 272 203 274 207
rect 274 203 277 207
rect 282 203 285 207
rect 285 203 287 207
rect 272 202 277 203
rect 282 202 287 203
rect 680 103 682 107
rect 682 103 685 107
rect 690 103 693 107
rect 693 103 695 107
rect 680 102 685 103
rect 690 102 695 103
rect 272 3 274 7
rect 274 3 277 7
rect 282 3 285 7
rect 285 3 287 7
rect 272 2 277 3
rect 282 2 287 3
<< metal6 >>
rect 272 807 288 830
rect 277 802 282 807
rect 287 802 288 807
rect 272 607 288 802
rect 277 602 282 607
rect 287 602 288 607
rect 272 407 288 602
rect 277 402 282 407
rect 287 402 288 407
rect 272 207 288 402
rect 277 202 282 207
rect 287 202 288 207
rect 272 7 288 202
rect 277 2 282 7
rect 287 2 288 7
rect 272 -30 288 2
rect 680 707 696 830
rect 685 702 690 707
rect 695 702 696 707
rect 680 507 696 702
rect 685 502 690 507
rect 695 502 696 507
rect 680 307 696 502
rect 685 302 690 307
rect 695 302 696 307
rect 680 107 696 302
rect 685 102 690 107
rect 695 102 696 107
rect 680 -30 696 102
use XOR2X1  XOR2X1_1
timestamp 1744883066
transform -1 0 60 0 -1 105
box -2 -3 58 103
use AND2X2  AND2X2_4
timestamp 1744883066
transform 1 0 60 0 -1 105
box -2 -3 34 103
use NOR3X1  NOR3X1_1
timestamp 1744883066
transform -1 0 68 0 1 105
box -2 -3 66 103
use OAI21X1  OAI21X1_5
timestamp 1744883066
transform 1 0 68 0 1 105
box -2 -3 34 103
use OR2X2  OR2X2_5
timestamp 1744883066
transform 1 0 92 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_1
timestamp 1744883066
transform -1 0 148 0 -1 105
box -2 -3 26 103
use NAND3X1  NAND3X1_1
timestamp 1744883066
transform -1 0 132 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_3
timestamp 1744883066
transform 1 0 132 0 1 105
box -2 -3 26 103
use AOI22X1  AOI22X1_8
timestamp 1744883066
transform 1 0 148 0 -1 105
box -2 -3 42 103
use NAND2X1  NAND2X1_7
timestamp 1744883066
transform -1 0 212 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_4
timestamp 1744883066
transform -1 0 180 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_2
timestamp 1744883066
transform 1 0 180 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_26
timestamp 1744883066
transform -1 0 236 0 -1 105
box -2 -3 26 103
use OAI22X1  OAI22X1_4
timestamp 1744883066
transform 1 0 236 0 -1 105
box -2 -3 42 103
use FILL  FILL_0_0_0
timestamp 1744883066
transform -1 0 284 0 -1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_3
timestamp 1744883066
transform -1 0 244 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_34
timestamp 1744883066
transform 1 0 244 0 1 105
box -2 -3 26 103
use FILL  FILL_1_0_0
timestamp 1744883066
transform 1 0 268 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_1
timestamp 1744883066
transform 1 0 276 0 1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1744883066
transform -1 0 292 0 -1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_27
timestamp 1744883066
transform -1 0 316 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_11
timestamp 1744883066
transform 1 0 316 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_6
timestamp 1744883066
transform -1 0 372 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_9
timestamp 1744883066
transform 1 0 284 0 1 105
box -2 -3 26 103
use NAND3X1  NAND3X1_3
timestamp 1744883066
transform 1 0 308 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_8
timestamp 1744883066
transform 1 0 340 0 1 105
box -2 -3 34 103
use OR2X2  OR2X2_1
timestamp 1744883066
transform -1 0 404 0 -1 105
box -2 -3 34 103
use AOI22X1  AOI22X1_4
timestamp 1744883066
transform 1 0 404 0 -1 105
box -2 -3 42 103
use NOR2X1  NOR2X1_5
timestamp 1744883066
transform 1 0 372 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_3
timestamp 1744883066
transform -1 0 428 0 1 105
box -2 -3 34 103
use AND2X2  AND2X2_5
timestamp 1744883066
transform -1 0 476 0 -1 105
box -2 -3 34 103
use XOR2X1  XOR2X1_3
timestamp 1744883066
transform 1 0 476 0 -1 105
box -2 -3 58 103
use AOI21X1  AOI21X1_4
timestamp 1744883066
transform 1 0 428 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_4
timestamp 1744883066
transform -1 0 492 0 1 105
box -2 -3 34 103
use BUFX2  BUFX2_6
timestamp 1744883066
transform 1 0 532 0 -1 105
box -2 -3 26 103
use AOI22X1  AOI22X1_5
timestamp 1744883066
transform -1 0 532 0 1 105
box -2 -3 42 103
use OAI21X1  OAI21X1_12
timestamp 1744883066
transform 1 0 532 0 1 105
box -2 -3 34 103
use BUFX2  BUFX2_3
timestamp 1744883066
transform 1 0 556 0 -1 105
box -2 -3 26 103
use XOR2X1  XOR2X1_4
timestamp 1744883066
transform -1 0 636 0 -1 105
box -2 -3 58 103
use NOR3X1  NOR3X1_4
timestamp 1744883066
transform 1 0 564 0 1 105
box -2 -3 66 103
use AOI22X1  AOI22X1_6
timestamp 1744883066
transform -1 0 676 0 -1 105
box -2 -3 42 103
use FILL  FILL_0_1_0
timestamp 1744883066
transform -1 0 684 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1744883066
transform -1 0 692 0 -1 105
box -2 -3 10 103
use NAND2X1  NAND2X1_11
timestamp 1744883066
transform -1 0 716 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_13
timestamp 1744883066
transform 1 0 628 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_16
timestamp 1744883066
transform -1 0 692 0 1 105
box -2 -3 34 103
use FILL  FILL_1_1_0
timestamp 1744883066
transform 1 0 692 0 1 105
box -2 -3 10 103
use INVX2  INVX2_8
timestamp 1744883066
transform 1 0 716 0 -1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_10
timestamp 1744883066
transform 1 0 732 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_4
timestamp 1744883066
transform 1 0 756 0 -1 105
box -2 -3 18 103
use FILL  FILL_1_1_1
timestamp 1744883066
transform 1 0 700 0 1 105
box -2 -3 10 103
use INVX2  INVX2_2
timestamp 1744883066
transform 1 0 708 0 1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_6
timestamp 1744883066
transform 1 0 724 0 1 105
box -2 -3 26 103
use INVX2  INVX2_3
timestamp 1744883066
transform -1 0 764 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_20
timestamp 1744883066
transform 1 0 772 0 -1 105
box -2 -3 34 103
use INVX2  INVX2_4
timestamp 1744883066
transform -1 0 820 0 -1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_19
timestamp 1744883066
transform 1 0 820 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_8
timestamp 1744883066
transform 1 0 764 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_25
timestamp 1744883066
transform -1 0 828 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_10
timestamp 1744883066
transform 1 0 828 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_8
timestamp 1744883066
transform -1 0 868 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_8
timestamp 1744883066
transform -1 0 892 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_6
timestamp 1744883066
transform -1 0 908 0 -1 105
box -2 -3 18 103
use AOI21X1  AOI21X1_5
timestamp 1744883066
transform -1 0 892 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_10
timestamp 1744883066
transform 1 0 892 0 1 105
box -2 -3 34 103
use XOR2X1  XOR2X1_2
timestamp 1744883066
transform -1 0 964 0 -1 105
box -2 -3 58 103
use FILL  FILL_1_1
timestamp 1744883066
transform -1 0 972 0 -1 105
box -2 -3 10 103
use AOI21X1  AOI21X1_10
timestamp 1744883066
transform -1 0 956 0 1 105
box -2 -3 34 103
use FILL  FILL_2_1
timestamp 1744883066
transform 1 0 956 0 1 105
box -2 -3 10 103
use FILL  FILL_2_2
timestamp 1744883066
transform 1 0 964 0 1 105
box -2 -3 10 103
use FILL  FILL_1_2
timestamp 1744883066
transform -1 0 980 0 -1 105
box -2 -3 10 103
use FILL  FILL_2_3
timestamp 1744883066
transform 1 0 972 0 1 105
box -2 -3 10 103
use BUFX2  BUFX2_5
timestamp 1744883066
transform -1 0 28 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_5
timestamp 1744883066
transform -1 0 52 0 -1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_9
timestamp 1744883066
transform -1 0 84 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_1
timestamp 1744883066
transform -1 0 116 0 -1 305
box -2 -3 34 103
use NOR3X1  NOR3X1_3
timestamp 1744883066
transform -1 0 180 0 -1 305
box -2 -3 66 103
use OAI21X1  OAI21X1_18
timestamp 1744883066
transform -1 0 212 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_6
timestamp 1744883066
transform -1 0 244 0 -1 305
box -2 -3 34 103
use OR2X2  OR2X2_2
timestamp 1744883066
transform 1 0 244 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_0_0
timestamp 1744883066
transform -1 0 284 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1744883066
transform -1 0 292 0 -1 305
box -2 -3 10 103
use NOR2X1  NOR2X1_1
timestamp 1744883066
transform -1 0 316 0 -1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_2
timestamp 1744883066
transform 1 0 316 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_45
timestamp 1744883066
transform 1 0 348 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_15
timestamp 1744883066
transform -1 0 396 0 -1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_24
timestamp 1744883066
transform 1 0 396 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_9
timestamp 1744883066
transform 1 0 420 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_14
timestamp 1744883066
transform -1 0 468 0 -1 305
box -2 -3 18 103
use AOI22X1  AOI22X1_3
timestamp 1744883066
transform 1 0 468 0 -1 305
box -2 -3 42 103
use INVX1  INVX1_1
timestamp 1744883066
transform 1 0 508 0 -1 305
box -2 -3 18 103
use AOI22X1  AOI22X1_7
timestamp 1744883066
transform -1 0 564 0 -1 305
box -2 -3 42 103
use AOI21X1  AOI21X1_15
timestamp 1744883066
transform 1 0 564 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_7
timestamp 1744883066
transform 1 0 596 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_14
timestamp 1744883066
transform 1 0 628 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_7
timestamp 1744883066
transform -1 0 684 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_1_0
timestamp 1744883066
transform -1 0 692 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1744883066
transform -1 0 700 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_15
timestamp 1744883066
transform -1 0 732 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_12
timestamp 1744883066
transform -1 0 756 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_29
timestamp 1744883066
transform -1 0 788 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_30
timestamp 1744883066
transform -1 0 812 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_9
timestamp 1744883066
transform 1 0 812 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_21
timestamp 1744883066
transform -1 0 876 0 -1 305
box -2 -3 34 103
use INVX2  INVX2_6
timestamp 1744883066
transform -1 0 892 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_13
timestamp 1744883066
transform -1 0 916 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_9
timestamp 1744883066
transform -1 0 940 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_19
timestamp 1744883066
transform -1 0 972 0 -1 305
box -2 -3 34 103
use FILL  FILL_3_1
timestamp 1744883066
transform -1 0 980 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_4
timestamp 1744883066
transform 1 0 4 0 1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_1
timestamp 1744883066
transform 1 0 36 0 1 305
box -2 -3 42 103
use INVX2  INVX2_12
timestamp 1744883066
transform 1 0 76 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_52
timestamp 1744883066
transform 1 0 92 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_3
timestamp 1744883066
transform 1 0 124 0 1 305
box -2 -3 26 103
use OR2X2  OR2X2_3
timestamp 1744883066
transform 1 0 148 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_1
timestamp 1744883066
transform 1 0 180 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_22
timestamp 1744883066
transform 1 0 212 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_4
timestamp 1744883066
transform -1 0 268 0 1 305
box -2 -3 26 103
use FILL  FILL_3_0_0
timestamp 1744883066
transform 1 0 268 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1744883066
transform 1 0 276 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_7
timestamp 1744883066
transform 1 0 284 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_8
timestamp 1744883066
transform -1 0 340 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_6
timestamp 1744883066
transform 1 0 340 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_31
timestamp 1744883066
transform 1 0 372 0 1 305
box -2 -3 34 103
use INVX1  INVX1_8
timestamp 1744883066
transform -1 0 420 0 1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_28
timestamp 1744883066
transform 1 0 420 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_27
timestamp 1744883066
transform 1 0 444 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_10
timestamp 1744883066
transform -1 0 500 0 1 305
box -2 -3 26 103
use AOI22X1  AOI22X1_9
timestamp 1744883066
transform 1 0 500 0 1 305
box -2 -3 42 103
use OAI21X1  OAI21X1_22
timestamp 1744883066
transform -1 0 572 0 1 305
box -2 -3 34 103
use INVX1  INVX1_2
timestamp 1744883066
transform -1 0 588 0 1 305
box -2 -3 18 103
use NOR3X1  NOR3X1_2
timestamp 1744883066
transform -1 0 652 0 1 305
box -2 -3 66 103
use OAI21X1  OAI21X1_24
timestamp 1744883066
transform 1 0 652 0 1 305
box -2 -3 34 103
use FILL  FILL_3_1_0
timestamp 1744883066
transform -1 0 692 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1744883066
transform -1 0 700 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_23
timestamp 1744883066
transform -1 0 732 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_14
timestamp 1744883066
transform -1 0 756 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_37
timestamp 1744883066
transform 1 0 756 0 1 305
box -2 -3 34 103
use INVX1  INVX1_7
timestamp 1744883066
transform 1 0 788 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_30
timestamp 1744883066
transform -1 0 836 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_36
timestamp 1744883066
transform -1 0 868 0 1 305
box -2 -3 34 103
use INVX2  INVX2_9
timestamp 1744883066
transform -1 0 884 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_42
timestamp 1744883066
transform 1 0 884 0 1 305
box -2 -3 34 103
use INVX1  INVX1_11
timestamp 1744883066
transform 1 0 916 0 1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_18
timestamp 1744883066
transform -1 0 956 0 1 305
box -2 -3 26 103
use FILL  FILL_4_1
timestamp 1744883066
transform 1 0 956 0 1 305
box -2 -3 10 103
use FILL  FILL_4_2
timestamp 1744883066
transform 1 0 964 0 1 305
box -2 -3 10 103
use FILL  FILL_4_3
timestamp 1744883066
transform 1 0 972 0 1 305
box -2 -3 10 103
use INVX2  INVX2_13
timestamp 1744883066
transform 1 0 4 0 -1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_26
timestamp 1744883066
transform 1 0 20 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_49
timestamp 1744883066
transform 1 0 44 0 -1 505
box -2 -3 34 103
use AND2X2  AND2X2_3
timestamp 1744883066
transform 1 0 76 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_25
timestamp 1744883066
transform -1 0 132 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_12
timestamp 1744883066
transform -1 0 164 0 -1 505
box -2 -3 34 103
use OR2X2  OR2X2_4
timestamp 1744883066
transform -1 0 196 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_2
timestamp 1744883066
transform 1 0 196 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_17
timestamp 1744883066
transform 1 0 228 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_31
timestamp 1744883066
transform -1 0 284 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_0_0
timestamp 1744883066
transform -1 0 292 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1744883066
transform -1 0 300 0 -1 505
box -2 -3 10 103
use NAND2X1  NAND2X1_32
timestamp 1744883066
transform -1 0 324 0 -1 505
box -2 -3 26 103
use AOI22X1  AOI22X1_2
timestamp 1744883066
transform -1 0 364 0 -1 505
box -2 -3 42 103
use NAND2X1  NAND2X1_33
timestamp 1744883066
transform 1 0 364 0 -1 505
box -2 -3 26 103
use AOI22X1  AOI22X1_12
timestamp 1744883066
transform -1 0 428 0 -1 505
box -2 -3 42 103
use OAI21X1  OAI21X1_47
timestamp 1744883066
transform -1 0 460 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_31
timestamp 1744883066
transform 1 0 460 0 -1 505
box -2 -3 26 103
use INVX2  INVX2_19
timestamp 1744883066
transform 1 0 484 0 -1 505
box -2 -3 18 103
use INVX2  INVX2_1
timestamp 1744883066
transform -1 0 516 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_33
timestamp 1744883066
transform -1 0 548 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_14
timestamp 1744883066
transform -1 0 580 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_14
timestamp 1744883066
transform 1 0 580 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_26
timestamp 1744883066
transform 1 0 612 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_28
timestamp 1744883066
transform 1 0 644 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_1_0
timestamp 1744883066
transform 1 0 676 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1744883066
transform 1 0 684 0 -1 505
box -2 -3 10 103
use AOI21X1  AOI21X1_11
timestamp 1744883066
transform 1 0 692 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_5
timestamp 1744883066
transform 1 0 724 0 -1 505
box -2 -3 34 103
use INVX2  INVX2_14
timestamp 1744883066
transform 1 0 756 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_32
timestamp 1744883066
transform 1 0 772 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_13
timestamp 1744883066
transform 1 0 804 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_12
timestamp 1744883066
transform 1 0 836 0 -1 505
box -2 -3 26 103
use NOR3X1  NOR3X1_5
timestamp 1744883066
transform -1 0 924 0 -1 505
box -2 -3 66 103
use BUFX2  BUFX2_9
timestamp 1744883066
transform 1 0 924 0 -1 505
box -2 -3 26 103
use AND2X2  AND2X2_2
timestamp 1744883066
transform 1 0 948 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_25
timestamp 1744883066
transform 1 0 4 0 1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_15
timestamp 1744883066
transform 1 0 28 0 1 505
box -2 -3 34 103
use AND2X2  AND2X2_6
timestamp 1744883066
transform 1 0 60 0 1 505
box -2 -3 34 103
use OAI22X1  OAI22X1_3
timestamp 1744883066
transform -1 0 132 0 1 505
box -2 -3 42 103
use NAND2X1  NAND2X1_21
timestamp 1744883066
transform 1 0 132 0 1 505
box -2 -3 26 103
use INVX2  INVX2_15
timestamp 1744883066
transform 1 0 156 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_50
timestamp 1744883066
transform 1 0 172 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_18
timestamp 1744883066
transform 1 0 204 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_51
timestamp 1744883066
transform -1 0 268 0 1 505
box -2 -3 34 103
use FILL  FILL_5_0_0
timestamp 1744883066
transform -1 0 276 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1744883066
transform -1 0 284 0 1 505
box -2 -3 10 103
use NOR2X1  NOR2X1_43
timestamp 1744883066
transform -1 0 308 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_30
timestamp 1744883066
transform -1 0 332 0 1 505
box -2 -3 26 103
use INVX1  INVX1_16
timestamp 1744883066
transform 1 0 332 0 1 505
box -2 -3 18 103
use AOI22X1  AOI22X1_11
timestamp 1744883066
transform 1 0 348 0 1 505
box -2 -3 42 103
use OAI21X1  OAI21X1_46
timestamp 1744883066
transform -1 0 420 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_39
timestamp 1744883066
transform -1 0 444 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_48
timestamp 1744883066
transform -1 0 476 0 1 505
box -2 -3 34 103
use INVX1  INVX1_3
timestamp 1744883066
transform 1 0 476 0 1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_15
timestamp 1744883066
transform -1 0 516 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_44
timestamp 1744883066
transform -1 0 548 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_43
timestamp 1744883066
transform -1 0 580 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_13
timestamp 1744883066
transform -1 0 604 0 1 505
box -2 -3 26 103
use OAI22X1  OAI22X1_1
timestamp 1744883066
transform -1 0 644 0 1 505
box -2 -3 42 103
use INVX1  INVX1_9
timestamp 1744883066
transform -1 0 660 0 1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_11
timestamp 1744883066
transform 1 0 660 0 1 505
box -2 -3 26 103
use FILL  FILL_5_1_0
timestamp 1744883066
transform -1 0 692 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1744883066
transform -1 0 700 0 1 505
box -2 -3 10 103
use NOR2X1  NOR2X1_29
timestamp 1744883066
transform -1 0 724 0 1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_8
timestamp 1744883066
transform 1 0 724 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_16
timestamp 1744883066
transform 1 0 756 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_23
timestamp 1744883066
transform 1 0 780 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_41
timestamp 1744883066
transform -1 0 836 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_22
timestamp 1744883066
transform -1 0 860 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_38
timestamp 1744883066
transform -1 0 892 0 1 505
box -2 -3 34 103
use INVX1  INVX1_13
timestamp 1744883066
transform -1 0 908 0 1 505
box -2 -3 18 103
use INVX2  INVX2_11
timestamp 1744883066
transform -1 0 924 0 1 505
box -2 -3 18 103
use BUFX2  BUFX2_11
timestamp 1744883066
transform 1 0 924 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_17
timestamp 1744883066
transform 1 0 948 0 1 505
box -2 -3 34 103
use NOR3X1  NOR3X1_8
timestamp 1744883066
transform -1 0 68 0 -1 705
box -2 -3 66 103
use NAND2X1  NAND2X1_27
timestamp 1744883066
transform -1 0 92 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_41
timestamp 1744883066
transform -1 0 116 0 -1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_16
timestamp 1744883066
transform -1 0 148 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_28
timestamp 1744883066
transform -1 0 172 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_29
timestamp 1744883066
transform -1 0 196 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_33
timestamp 1744883066
transform 1 0 196 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_36
timestamp 1744883066
transform -1 0 244 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_37
timestamp 1744883066
transform 1 0 244 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_0_0
timestamp 1744883066
transform 1 0 268 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1744883066
transform 1 0 276 0 -1 705
box -2 -3 10 103
use NOR2X1  NOR2X1_40
timestamp 1744883066
transform 1 0 284 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_38
timestamp 1744883066
transform 1 0 308 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_42
timestamp 1744883066
transform 1 0 332 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_34
timestamp 1744883066
transform 1 0 356 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_44
timestamp 1744883066
transform -1 0 404 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_35
timestamp 1744883066
transform 1 0 404 0 -1 705
box -2 -3 26 103
use INVX2  INVX2_17
timestamp 1744883066
transform 1 0 428 0 -1 705
box -2 -3 18 103
use AOI22X1  AOI22X1_10
timestamp 1744883066
transform -1 0 484 0 -1 705
box -2 -3 42 103
use OAI21X1  OAI21X1_39
timestamp 1744883066
transform -1 0 516 0 -1 705
box -2 -3 34 103
use INVX2  INVX2_5
timestamp 1744883066
transform 1 0 516 0 -1 705
box -2 -3 18 103
use AOI21X1  AOI21X1_21
timestamp 1744883066
transform -1 0 564 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_34
timestamp 1744883066
transform -1 0 596 0 -1 705
box -2 -3 34 103
use OAI22X1  OAI22X1_2
timestamp 1744883066
transform 1 0 596 0 -1 705
box -2 -3 42 103
use NOR2X1  NOR2X1_15
timestamp 1744883066
transform 1 0 636 0 -1 705
box -2 -3 26 103
use INVX2  INVX2_7
timestamp 1744883066
transform 1 0 660 0 -1 705
box -2 -3 18 103
use FILL  FILL_6_1_0
timestamp 1744883066
transform 1 0 676 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1744883066
transform 1 0 684 0 -1 705
box -2 -3 10 103
use NAND3X1  NAND3X1_12
timestamp 1744883066
transform 1 0 692 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_16
timestamp 1744883066
transform 1 0 724 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_35
timestamp 1744883066
transform 1 0 748 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_21
timestamp 1744883066
transform 1 0 780 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_14
timestamp 1744883066
transform 1 0 804 0 -1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_7
timestamp 1744883066
transform -1 0 860 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_16
timestamp 1744883066
transform -1 0 892 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_19
timestamp 1744883066
transform -1 0 924 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_5
timestamp 1744883066
transform -1 0 940 0 -1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_17
timestamp 1744883066
transform -1 0 964 0 -1 705
box -2 -3 26 103
use FILL  FILL_7_1
timestamp 1744883066
transform -1 0 972 0 -1 705
box -2 -3 10 103
use FILL  FILL_7_2
timestamp 1744883066
transform -1 0 980 0 -1 705
box -2 -3 10 103
use BUFX2  BUFX2_4
timestamp 1744883066
transform -1 0 28 0 1 705
box -2 -3 26 103
use INVX1  INVX1_20
timestamp 1744883066
transform -1 0 44 0 1 705
box -2 -3 18 103
use INVX1  INVX1_18
timestamp 1744883066
transform 1 0 44 0 1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_23
timestamp 1744883066
transform -1 0 84 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_20
timestamp 1744883066
transform 1 0 84 0 1 705
box -2 -3 26 103
use INVX1  INVX1_17
timestamp 1744883066
transform 1 0 108 0 1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_17
timestamp 1744883066
transform -1 0 148 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_22
timestamp 1744883066
transform 1 0 148 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_2
timestamp 1744883066
transform 1 0 172 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_2
timestamp 1744883066
transform 1 0 196 0 1 705
box -2 -3 26 103
use AND2X2  AND2X2_1
timestamp 1744883066
transform -1 0 252 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_24
timestamp 1744883066
transform 1 0 252 0 1 705
box -2 -3 26 103
use FILL  FILL_7_0_0
timestamp 1744883066
transform -1 0 284 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1744883066
transform -1 0 292 0 1 705
box -2 -3 10 103
use INVX1  INVX1_19
timestamp 1744883066
transform -1 0 308 0 1 705
box -2 -3 18 103
use INVX2  INVX2_16
timestamp 1744883066
transform -1 0 324 0 1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_32
timestamp 1744883066
transform -1 0 348 0 1 705
box -2 -3 26 103
use INVX2  INVX2_18
timestamp 1744883066
transform -1 0 364 0 1 705
box -2 -3 18 103
use NAND3X1  NAND3X1_13
timestamp 1744883066
transform 1 0 364 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_20
timestamp 1744883066
transform -1 0 428 0 1 705
box -2 -3 34 103
use INVX1  INVX1_12
timestamp 1744883066
transform -1 0 444 0 1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_18
timestamp 1744883066
transform 1 0 444 0 1 705
box -2 -3 26 103
use INVX2  INVX2_10
timestamp 1744883066
transform -1 0 484 0 1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_19
timestamp 1744883066
transform 1 0 484 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_20
timestamp 1744883066
transform -1 0 532 0 1 705
box -2 -3 26 103
use INVX4  INVX4_1
timestamp 1744883066
transform 1 0 532 0 1 705
box -2 -3 26 103
use NOR3X1  NOR3X1_6
timestamp 1744883066
transform -1 0 620 0 1 705
box -2 -3 66 103
use AOI21X1  AOI21X1_17
timestamp 1744883066
transform -1 0 652 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_40
timestamp 1744883066
transform -1 0 684 0 1 705
box -2 -3 34 103
use FILL  FILL_7_1_0
timestamp 1744883066
transform 1 0 684 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1744883066
transform 1 0 692 0 1 705
box -2 -3 10 103
use NAND3X1  NAND3X1_11
timestamp 1744883066
transform 1 0 700 0 1 705
box -2 -3 34 103
use INVX1  INVX1_10
timestamp 1744883066
transform -1 0 748 0 1 705
box -2 -3 18 103
use NAND3X1  NAND3X1_6
timestamp 1744883066
transform -1 0 780 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_18
timestamp 1744883066
transform 1 0 780 0 1 705
box -2 -3 34 103
use NOR3X1  NOR3X1_7
timestamp 1744883066
transform 1 0 812 0 1 705
box -2 -3 66 103
use BUFX2  BUFX2_2
timestamp 1744883066
transform 1 0 876 0 1 705
box -2 -3 26 103
use BUFX2  BUFX2_1
timestamp 1744883066
transform 1 0 900 0 1 705
box -2 -3 26 103
use BUFX2  BUFX2_7
timestamp 1744883066
transform 1 0 924 0 1 705
box -2 -3 26 103
use BUFX2  BUFX2_10
timestamp 1744883066
transform -1 0 972 0 1 705
box -2 -3 26 103
use FILL  FILL_8_1
timestamp 1744883066
transform 1 0 972 0 1 705
box -2 -3 10 103
<< labels >>
flabel metal6 s 272 -30 288 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 680 -30 696 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal3 s -26 568 -22 572 7 FreeSans 24 0 0 0 A[0]
port 2 nsew
flabel metal3 s -26 468 -22 472 7 FreeSans 24 0 0 0 A[1]
port 3 nsew
flabel metal3 s -26 88 -22 92 7 FreeSans 24 0 0 0 A[2]
port 4 nsew
flabel metal2 s 334 -22 338 -18 7 FreeSans 24 270 0 0 A[3]
port 5 nsew
flabel metal2 s 734 -22 738 -18 7 FreeSans 24 270 0 0 A[4]
port 6 nsew
flabel metal3 s 1006 338 1010 342 3 FreeSans 24 0 0 0 A[5]
port 7 nsew
flabel metal3 s 1006 578 1010 582 3 FreeSans 24 0 0 0 A[6]
port 8 nsew
flabel metal2 s 494 828 498 832 3 FreeSans 24 90 0 0 A[7]
port 9 nsew
flabel metal3 s -26 548 -22 552 7 FreeSans 24 0 0 0 B[0]
port 10 nsew
flabel metal3 s -26 448 -22 452 7 FreeSans 24 0 0 0 B[1]
port 11 nsew
flabel metal3 s -26 68 -22 72 7 FreeSans 24 0 0 0 B[2]
port 12 nsew
flabel metal2 s 470 -22 474 -18 7 FreeSans 24 270 0 0 B[3]
port 13 nsew
flabel metal2 s 630 -22 634 -18 7 FreeSans 24 270 0 0 B[4]
port 14 nsew
flabel metal3 s 1006 258 1010 262 3 FreeSans 24 0 0 0 B[5]
port 15 nsew
flabel metal3 s 1006 558 1010 562 3 FreeSans 24 0 0 0 B[6]
port 16 nsew
flabel metal2 s 470 828 474 832 3 FreeSans 24 90 0 0 B[7]
port 17 nsew
flabel metal3 s -26 738 -22 742 7 FreeSans 24 90 0 0 opcode[0]
port 18 nsew
flabel metal2 s 102 828 106 832 3 FreeSans 24 90 0 0 opcode[1]
port 19 nsew
flabel metal2 s 326 828 330 832 3 FreeSans 24 90 0 0 opcode[2]
port 20 nsew
flabel metal2 s 350 828 354 832 3 FreeSans 24 90 0 0 opcode[3]
port 21 nsew
flabel metal2 s 566 -22 570 -18 7 FreeSans 24 270 0 0 result[0]
port 22 nsew
flabel metal3 s -26 758 -22 762 7 FreeSans 24 90 0 0 result[1]
port 23 nsew
flabel metal3 s -26 248 -22 252 7 FreeSans 24 0 0 0 result[2]
port 24 nsew
flabel metal2 s 542 -22 546 -18 7 FreeSans 24 270 0 0 result[3]
port 25 nsew
flabel metal2 s 934 -22 938 -18 3 FreeSans 24 270 0 0 result[4]
port 26 nsew
flabel metal2 s 878 -22 882 -18 7 FreeSans 24 270 0 0 result[5]
port 27 nsew
flabel metal3 s 1006 448 1010 452 3 FreeSans 24 0 0 0 result[6]
port 28 nsew
flabel metal2 s 958 828 962 832 3 FreeSans 24 90 0 0 result[7]
port 29 nsew
flabel metal2 s 886 828 890 832 3 FreeSans 24 90 0 0 overflow
port 30 nsew
flabel metal2 s 910 828 914 832 3 FreeSans 24 90 0 0 negative
port 31 nsew
flabel metal3 s 1006 598 1010 602 3 FreeSans 24 0 0 0 zero
port 32 nsew
<< end >>
