magic
tech scmos
timestamp 1743078376
<< metal1 >>
rect 608 703 610 707
rect 614 703 617 707
rect 621 703 624 707
rect 306 678 321 681
rect 634 678 641 681
rect 38 671 41 678
rect 26 668 33 671
rect 38 668 49 671
rect 54 668 70 671
rect 150 671 153 678
rect 318 672 321 678
rect 150 668 161 671
rect 214 668 222 671
rect 350 668 361 671
rect 394 668 401 671
rect 518 668 545 671
rect 582 668 590 671
rect 646 668 657 671
rect 806 668 817 671
rect 806 662 809 668
rect 94 658 110 661
rect 182 658 201 661
rect 362 658 369 661
rect 442 658 449 661
rect 554 658 561 661
rect 594 658 601 661
rect 22 648 33 651
rect 182 648 185 658
rect 294 651 297 658
rect 286 648 297 651
rect 830 648 841 651
rect 114 638 115 642
rect 141 618 142 622
rect 238 618 254 621
rect 602 618 603 622
rect 232 603 234 607
rect 238 603 241 607
rect 245 603 248 607
rect 733 588 734 592
rect 870 581 873 588
rect 862 578 873 581
rect 14 548 22 551
rect 46 551 49 561
rect 134 558 145 561
rect 150 558 169 561
rect 390 558 401 561
rect 430 558 438 561
rect 526 561 529 568
rect 830 562 834 564
rect 518 558 529 561
rect 42 548 49 551
rect 250 548 257 551
rect 326 548 337 551
rect 382 548 393 551
rect 482 548 489 551
rect 542 551 545 558
rect 814 552 818 554
rect 530 548 537 551
rect 542 548 553 551
rect 558 548 577 551
rect 142 541 145 548
rect 326 542 329 548
rect 390 542 393 548
rect 118 538 137 541
rect 142 538 153 541
rect 214 538 230 541
rect 242 538 249 541
rect 398 538 417 541
rect 574 538 577 548
rect 662 542 665 551
rect 694 548 702 551
rect 686 538 694 541
rect 766 538 774 541
rect 822 538 834 541
rect 22 528 25 538
rect 118 528 121 538
rect 566 528 569 538
rect 822 532 825 538
rect 652 528 654 532
rect 53 518 54 522
rect 298 518 300 522
rect 426 518 427 522
rect 622 521 625 528
rect 606 518 625 521
rect 608 503 610 507
rect 614 503 617 507
rect 621 503 624 507
rect 278 478 289 481
rect 470 478 486 481
rect 506 478 513 481
rect 218 468 225 471
rect 286 468 297 471
rect 598 468 625 471
rect 670 468 686 471
rect 838 468 854 471
rect 286 462 289 468
rect 598 462 601 468
rect 66 458 73 461
rect 78 458 105 461
rect 214 458 265 461
rect 314 458 321 461
rect 338 458 345 461
rect 426 458 433 461
rect 446 458 462 461
rect 482 458 489 461
rect 182 448 193 451
rect 322 448 326 452
rect 430 448 433 458
rect 726 451 729 458
rect 718 448 729 451
rect 590 438 622 441
rect 418 428 419 432
rect 232 403 234 407
rect 238 403 241 407
rect 245 403 248 407
rect 602 388 603 392
rect 557 368 558 372
rect 766 371 769 381
rect 766 368 785 371
rect 826 368 827 372
rect 38 348 62 351
rect 142 351 145 361
rect 250 358 257 361
rect 398 358 409 361
rect 614 358 630 361
rect 782 358 785 368
rect 406 352 409 358
rect 122 348 129 351
rect 142 348 161 351
rect 170 348 185 351
rect 278 348 286 351
rect 330 348 337 351
rect 210 338 217 341
rect 374 341 377 351
rect 454 351 457 358
rect 414 348 441 351
rect 454 348 465 351
rect 486 342 489 351
rect 506 348 513 351
rect 534 348 542 351
rect 678 348 686 351
rect 698 348 705 351
rect 734 348 745 351
rect 742 342 745 348
rect 362 338 377 341
rect 626 338 641 341
rect 690 338 697 341
rect 804 338 806 342
rect 862 338 870 341
rect 286 331 289 338
rect 286 328 297 331
rect 486 328 497 331
rect 670 331 673 338
rect 662 328 673 331
rect 317 318 318 322
rect 346 318 347 322
rect 608 303 610 307
rect 614 303 617 307
rect 621 303 624 307
rect 69 288 70 292
rect 306 278 313 281
rect 602 278 625 281
rect 782 278 790 281
rect 158 268 177 271
rect 406 268 425 271
rect 526 268 537 271
rect 690 268 705 271
rect 134 258 150 261
rect 230 258 265 261
rect 270 258 286 261
rect 302 258 313 261
rect 422 258 425 268
rect 558 258 566 261
rect 582 258 614 261
rect 678 258 694 261
rect 750 258 761 261
rect 230 248 233 258
rect 854 248 862 251
rect 510 238 518 241
rect 36 218 38 222
rect 186 218 187 222
rect 218 218 219 222
rect 298 218 299 222
rect 466 218 467 222
rect 557 218 558 222
rect 232 203 234 207
rect 238 203 241 207
rect 245 203 248 207
rect 573 168 574 172
rect 74 158 78 162
rect 86 158 97 161
rect 330 158 334 162
rect 830 161 833 168
rect 830 158 841 161
rect 22 148 33 151
rect 66 148 73 151
rect 118 148 126 151
rect 250 148 265 151
rect 574 148 582 151
rect 634 148 649 151
rect 802 148 809 151
rect 126 138 129 148
rect 358 138 377 141
rect 390 138 393 148
rect 454 138 465 141
rect 358 132 361 138
rect 454 132 457 138
rect 614 118 630 121
rect 608 103 610 107
rect 614 103 617 107
rect 621 103 624 107
rect 180 88 182 92
rect 236 88 238 92
rect 290 88 291 92
rect 557 88 558 92
rect 716 88 718 92
rect 458 78 462 82
rect 602 78 617 81
rect 622 78 641 81
rect 198 68 209 71
rect 398 68 409 71
rect 502 68 510 71
rect 566 68 574 71
rect 582 68 606 71
rect 678 68 689 71
rect 206 62 209 68
rect 62 58 97 61
rect 102 58 110 61
rect 294 58 313 61
rect 366 58 385 61
rect 414 61 417 68
rect 414 58 433 61
rect 526 61 529 68
rect 526 58 537 61
rect 774 58 790 61
rect 806 58 825 61
rect 830 58 849 61
rect 110 48 121 51
rect 294 48 297 58
rect 462 48 481 51
rect 526 48 537 51
rect 546 48 553 51
rect 642 48 649 51
rect 550 42 554 44
rect 232 3 234 7
rect 238 3 241 7
rect 245 3 248 7
<< m2contact >>
rect 610 703 614 707
rect 617 703 621 707
rect 486 688 490 692
rect 782 688 786 692
rect 38 678 42 682
rect 86 678 90 682
rect 150 678 154 682
rect 222 678 226 682
rect 334 678 338 682
rect 390 678 394 682
rect 550 678 554 682
rect 630 678 634 682
rect 790 678 794 682
rect 846 678 850 682
rect 6 668 10 672
rect 22 668 26 672
rect 70 668 74 672
rect 102 668 106 672
rect 182 668 186 672
rect 222 668 226 672
rect 262 668 266 672
rect 294 668 298 672
rect 318 668 322 672
rect 342 668 346 672
rect 374 668 378 672
rect 390 668 394 672
rect 422 668 426 672
rect 430 668 434 672
rect 462 668 466 672
rect 502 668 506 672
rect 590 668 594 672
rect 670 668 674 672
rect 686 668 690 672
rect 734 668 738 672
rect 758 668 762 672
rect 110 658 114 662
rect 134 658 138 662
rect 166 658 170 662
rect 206 658 210 662
rect 238 658 242 662
rect 270 658 274 662
rect 294 658 298 662
rect 318 658 322 662
rect 358 658 362 662
rect 438 658 442 662
rect 454 658 458 662
rect 470 658 474 662
rect 494 658 498 662
rect 526 658 530 662
rect 534 658 538 662
rect 550 658 554 662
rect 574 658 578 662
rect 590 658 594 662
rect 662 658 666 662
rect 806 658 810 662
rect 62 648 66 652
rect 126 648 130 652
rect 190 648 194 652
rect 310 648 314 652
rect 382 648 386 652
rect 414 648 418 652
rect 438 648 442 652
rect 678 648 682 652
rect 742 648 746 652
rect 750 648 754 652
rect 110 638 114 642
rect 614 638 618 642
rect 14 618 18 622
rect 78 618 82 622
rect 142 618 146 622
rect 254 618 258 622
rect 350 618 354 622
rect 430 618 434 622
rect 558 618 562 622
rect 598 618 602 622
rect 710 618 714 622
rect 806 618 810 622
rect 822 618 826 622
rect 234 603 238 607
rect 241 603 245 607
rect 342 588 346 592
rect 734 588 738 592
rect 870 588 874 592
rect 526 568 530 572
rect 582 568 586 572
rect 646 568 650 572
rect 22 548 26 552
rect 38 548 42 552
rect 270 558 274 562
rect 438 558 442 562
rect 454 558 458 562
rect 542 558 546 562
rect 606 558 610 562
rect 630 558 634 562
rect 718 558 722 562
rect 830 558 834 562
rect 94 548 98 552
rect 102 548 106 552
rect 142 548 146 552
rect 182 548 186 552
rect 222 548 226 552
rect 246 548 250 552
rect 366 548 370 552
rect 478 548 482 552
rect 526 548 530 552
rect 638 548 642 552
rect 6 538 10 542
rect 22 538 26 542
rect 62 538 66 542
rect 86 538 90 542
rect 158 538 162 542
rect 190 538 194 542
rect 230 538 234 542
rect 238 538 242 542
rect 262 538 266 542
rect 278 538 282 542
rect 326 538 330 542
rect 342 538 346 542
rect 358 538 362 542
rect 374 538 378 542
rect 390 538 394 542
rect 438 538 442 542
rect 510 538 514 542
rect 526 538 530 542
rect 566 538 570 542
rect 678 548 682 552
rect 702 548 706 552
rect 734 548 738 552
rect 750 548 754 552
rect 806 548 810 552
rect 814 548 818 552
rect 822 548 826 552
rect 846 548 850 552
rect 590 538 594 542
rect 662 538 666 542
rect 670 538 674 542
rect 694 538 698 542
rect 710 538 714 542
rect 742 538 746 542
rect 758 538 762 542
rect 774 538 778 542
rect 798 538 802 542
rect 70 528 74 532
rect 126 528 130 532
rect 198 528 202 532
rect 406 528 410 532
rect 462 528 466 532
rect 502 528 506 532
rect 622 528 626 532
rect 654 528 658 532
rect 774 528 778 532
rect 782 528 786 532
rect 822 528 826 532
rect 30 518 34 522
rect 54 518 58 522
rect 78 518 82 522
rect 110 518 114 522
rect 166 518 170 522
rect 206 518 210 522
rect 294 518 298 522
rect 422 518 426 522
rect 454 518 458 522
rect 470 518 474 522
rect 494 518 498 522
rect 790 518 794 522
rect 610 503 614 507
rect 617 503 621 507
rect 126 488 130 492
rect 430 488 434 492
rect 638 488 642 492
rect 814 488 818 492
rect 854 488 858 492
rect 30 478 34 482
rect 190 478 194 482
rect 406 478 410 482
rect 462 478 466 482
rect 486 478 490 482
rect 502 478 506 482
rect 518 478 522 482
rect 774 478 778 482
rect 822 478 826 482
rect 46 468 50 472
rect 86 468 90 472
rect 118 468 122 472
rect 150 468 154 472
rect 158 468 162 472
rect 174 468 178 472
rect 206 468 210 472
rect 214 468 218 472
rect 230 468 234 472
rect 254 468 258 472
rect 310 468 314 472
rect 350 468 354 472
rect 366 468 370 472
rect 398 468 402 472
rect 454 468 458 472
rect 558 468 562 472
rect 574 468 578 472
rect 654 468 658 472
rect 686 468 690 472
rect 702 468 706 472
rect 726 468 730 472
rect 798 468 802 472
rect 854 468 858 472
rect 870 468 874 472
rect 22 458 26 462
rect 38 458 42 462
rect 54 458 58 462
rect 62 458 66 462
rect 110 458 114 462
rect 142 458 146 462
rect 166 458 170 462
rect 286 458 290 462
rect 302 458 306 462
rect 310 458 314 462
rect 334 458 338 462
rect 374 458 378 462
rect 422 458 426 462
rect 462 458 466 462
rect 478 458 482 462
rect 494 458 498 462
rect 526 458 530 462
rect 542 458 546 462
rect 550 458 554 462
rect 598 458 602 462
rect 646 458 650 462
rect 662 458 666 462
rect 678 458 682 462
rect 726 458 730 462
rect 750 458 754 462
rect 782 458 786 462
rect 846 458 850 462
rect 62 448 66 452
rect 94 448 98 452
rect 278 448 282 452
rect 318 448 322 452
rect 334 448 338 452
rect 350 448 354 452
rect 390 448 394 452
rect 534 448 538 452
rect 582 448 586 452
rect 638 448 642 452
rect 710 448 714 452
rect 758 448 762 452
rect 790 448 794 452
rect 814 448 818 452
rect 854 448 858 452
rect 6 438 10 442
rect 622 438 626 442
rect 742 438 746 442
rect 774 438 778 442
rect 414 428 418 432
rect 750 428 754 432
rect 478 418 482 422
rect 566 418 570 422
rect 694 418 698 422
rect 822 418 826 422
rect 234 403 238 407
rect 241 403 245 407
rect 598 388 602 392
rect 558 368 562 372
rect 758 368 762 372
rect 798 368 802 372
rect 822 368 826 372
rect 62 358 66 362
rect 110 358 114 362
rect 62 348 66 352
rect 78 348 82 352
rect 118 348 122 352
rect 198 358 202 362
rect 246 358 250 362
rect 310 358 314 362
rect 422 358 426 362
rect 454 358 458 362
rect 542 358 546 362
rect 630 358 634 362
rect 662 358 666 362
rect 718 358 722 362
rect 742 358 746 362
rect 774 358 778 362
rect 838 358 842 362
rect 166 348 170 352
rect 206 348 210 352
rect 286 348 290 352
rect 326 348 330 352
rect 366 348 370 352
rect 6 338 10 342
rect 54 338 58 342
rect 86 338 90 342
rect 94 338 98 342
rect 118 338 122 342
rect 174 338 178 342
rect 206 338 210 342
rect 286 338 290 342
rect 326 338 330 342
rect 342 338 346 342
rect 358 338 362 342
rect 406 348 410 352
rect 502 348 506 352
rect 542 348 546 352
rect 558 348 562 352
rect 598 348 602 352
rect 646 348 650 352
rect 670 348 674 352
rect 686 348 690 352
rect 694 348 698 352
rect 710 348 714 352
rect 766 348 770 352
rect 790 348 794 352
rect 822 348 826 352
rect 846 348 850 352
rect 382 338 386 342
rect 406 338 410 342
rect 430 338 434 342
rect 470 338 474 342
rect 486 338 490 342
rect 518 338 522 342
rect 566 338 570 342
rect 574 338 578 342
rect 590 338 594 342
rect 622 338 626 342
rect 670 338 674 342
rect 686 338 690 342
rect 726 338 730 342
rect 742 338 746 342
rect 806 338 810 342
rect 814 338 818 342
rect 870 338 874 342
rect 150 328 154 332
rect 230 328 234 332
rect 262 328 266 332
rect 270 328 274 332
rect 302 328 306 332
rect 398 328 402 332
rect 454 328 458 332
rect 502 328 506 332
rect 534 328 538 332
rect 686 328 690 332
rect 62 318 66 322
rect 110 318 114 322
rect 142 318 146 322
rect 198 318 202 322
rect 222 318 226 322
rect 318 318 322 322
rect 342 318 346 322
rect 582 318 586 322
rect 610 303 614 307
rect 617 303 621 307
rect 70 288 74 292
rect 350 288 354 292
rect 726 288 730 292
rect 774 288 778 292
rect 150 278 154 282
rect 286 278 290 282
rect 302 278 306 282
rect 398 278 402 282
rect 446 278 450 282
rect 510 278 514 282
rect 518 278 522 282
rect 598 278 602 282
rect 630 278 634 282
rect 742 278 746 282
rect 790 278 794 282
rect 6 268 10 272
rect 54 268 58 272
rect 78 268 82 272
rect 118 268 122 272
rect 206 268 210 272
rect 278 268 282 272
rect 318 268 322 272
rect 326 268 330 272
rect 366 268 370 272
rect 382 268 386 272
rect 430 268 434 272
rect 454 268 458 272
rect 494 268 498 272
rect 566 268 570 272
rect 574 268 578 272
rect 638 268 642 272
rect 654 268 658 272
rect 686 268 690 272
rect 710 268 714 272
rect 734 268 738 272
rect 766 268 770 272
rect 806 268 810 272
rect 822 268 826 272
rect 838 268 842 272
rect 102 258 106 262
rect 126 258 130 262
rect 150 258 154 262
rect 166 258 170 262
rect 182 258 186 262
rect 214 258 218 262
rect 286 258 290 262
rect 334 258 338 262
rect 358 258 362 262
rect 390 258 394 262
rect 414 258 418 262
rect 462 258 466 262
rect 486 258 490 262
rect 542 258 546 262
rect 566 258 570 262
rect 614 258 618 262
rect 646 258 650 262
rect 694 258 698 262
rect 814 258 818 262
rect 62 248 66 252
rect 86 248 90 252
rect 142 248 146 252
rect 198 248 202 252
rect 254 248 258 252
rect 350 248 354 252
rect 478 248 482 252
rect 590 248 594 252
rect 662 248 666 252
rect 670 248 674 252
rect 694 248 698 252
rect 798 248 802 252
rect 830 248 834 252
rect 862 248 866 252
rect 102 238 106 242
rect 518 238 522 242
rect 38 218 42 222
rect 94 218 98 222
rect 182 218 186 222
rect 214 218 218 222
rect 294 218 298 222
rect 366 218 370 222
rect 446 218 450 222
rect 462 218 466 222
rect 526 218 530 222
rect 558 218 562 222
rect 846 218 850 222
rect 234 203 238 207
rect 241 203 245 207
rect 310 188 314 192
rect 350 188 354 192
rect 854 188 858 192
rect 38 168 42 172
rect 574 168 578 172
rect 830 168 834 172
rect 54 158 58 162
rect 70 158 74 162
rect 150 158 154 162
rect 206 158 210 162
rect 222 158 226 162
rect 254 158 258 162
rect 326 158 330 162
rect 342 158 346 162
rect 390 158 394 162
rect 558 158 562 162
rect 662 158 666 162
rect 798 158 802 162
rect 46 148 50 152
rect 62 148 66 152
rect 126 148 130 152
rect 134 148 138 152
rect 158 148 162 152
rect 190 148 194 152
rect 230 148 234 152
rect 246 148 250 152
rect 270 148 274 152
rect 286 148 290 152
rect 326 148 330 152
rect 382 148 386 152
rect 390 148 394 152
rect 406 148 410 152
rect 454 148 458 152
rect 486 148 490 152
rect 502 148 506 152
rect 518 148 522 152
rect 534 148 538 152
rect 550 148 554 152
rect 582 148 586 152
rect 630 148 634 152
rect 670 148 674 152
rect 686 148 690 152
rect 702 148 706 152
rect 742 148 746 152
rect 782 148 786 152
rect 790 148 794 152
rect 798 148 802 152
rect 822 148 826 152
rect 6 138 10 142
rect 62 138 66 142
rect 110 138 114 142
rect 182 138 186 142
rect 198 138 202 142
rect 278 138 282 142
rect 294 138 298 142
rect 318 138 322 142
rect 414 138 418 142
rect 438 140 442 144
rect 446 138 450 142
rect 478 138 482 142
rect 494 138 498 142
rect 510 138 514 142
rect 526 138 530 142
rect 542 138 546 142
rect 582 138 586 142
rect 590 138 594 142
rect 598 140 602 144
rect 638 138 642 142
rect 678 138 682 142
rect 694 138 698 142
rect 718 138 722 142
rect 750 138 754 142
rect 774 138 778 142
rect 830 138 834 142
rect 862 138 866 142
rect 94 128 98 132
rect 174 128 178 132
rect 214 128 218 132
rect 310 128 314 132
rect 358 128 362 132
rect 366 128 370 132
rect 454 128 458 132
rect 470 128 474 132
rect 710 128 714 132
rect 766 128 770 132
rect 846 128 850 132
rect 150 118 154 122
rect 166 118 170 122
rect 422 118 426 122
rect 630 118 634 122
rect 662 118 666 122
rect 734 118 738 122
rect 758 118 762 122
rect 610 103 614 107
rect 617 103 621 107
rect 182 88 186 92
rect 238 88 242 92
rect 286 88 290 92
rect 310 88 314 92
rect 342 88 346 92
rect 526 88 530 92
rect 558 88 562 92
rect 718 88 722 92
rect 414 78 418 82
rect 454 78 458 82
rect 542 78 546 82
rect 598 78 602 82
rect 798 78 802 82
rect 30 68 34 72
rect 78 68 82 72
rect 86 68 90 72
rect 134 66 138 70
rect 142 68 146 72
rect 254 68 258 72
rect 278 68 282 72
rect 302 68 306 72
rect 318 68 322 72
rect 414 68 418 72
rect 446 68 450 72
rect 470 68 474 72
rect 486 68 490 72
rect 510 68 514 72
rect 526 68 530 72
rect 574 68 578 72
rect 606 68 610 72
rect 654 68 658 72
rect 734 68 738 72
rect 742 68 746 72
rect 790 68 794 72
rect 814 68 818 72
rect 22 58 26 62
rect 110 58 114 62
rect 206 58 210 62
rect 326 58 330 62
rect 390 58 394 62
rect 438 58 442 62
rect 494 58 498 62
rect 630 58 634 62
rect 662 58 666 62
rect 790 58 794 62
rect 374 48 378 52
rect 422 48 426 52
rect 454 48 458 52
rect 542 48 546 52
rect 638 48 642 52
rect 678 48 682 52
rect 838 48 842 52
rect 6 38 10 42
rect 550 38 554 42
rect 350 18 354 22
rect 862 18 866 22
rect 234 3 238 7
rect 241 3 245 7
<< metal2 >>
rect 150 728 154 732
rect 222 728 226 732
rect 302 728 306 732
rect 326 728 330 732
rect 478 731 482 732
rect 510 731 514 732
rect 478 728 489 731
rect 510 728 521 731
rect 150 702 153 728
rect 38 682 41 698
rect 150 682 153 698
rect 222 682 225 728
rect 302 692 305 728
rect 326 702 329 728
rect 294 688 302 691
rect 26 668 30 671
rect 6 652 9 668
rect 58 648 62 651
rect 14 562 17 618
rect 18 548 22 551
rect 34 548 38 551
rect 6 542 9 548
rect 6 522 9 538
rect 22 532 25 538
rect 30 482 33 518
rect 46 492 49 558
rect 54 522 57 538
rect 62 532 65 538
rect 70 532 73 668
rect 86 652 89 678
rect 98 668 102 671
rect 106 658 110 661
rect 130 658 134 661
rect 110 632 113 638
rect 78 572 81 618
rect 126 582 129 648
rect 142 562 145 618
rect 150 592 153 678
rect 178 668 182 671
rect 206 662 209 678
rect 222 672 225 678
rect 166 652 169 658
rect 190 642 193 648
rect 222 632 225 668
rect 238 662 241 678
rect 294 672 297 688
rect 318 672 321 678
rect 334 672 337 678
rect 342 672 345 698
rect 486 692 489 728
rect 258 668 262 671
rect 314 658 318 661
rect 254 622 257 658
rect 270 622 273 658
rect 294 652 297 658
rect 310 642 313 648
rect 342 642 345 668
rect 358 662 361 688
rect 386 678 390 681
rect 382 668 390 671
rect 374 662 377 668
rect 382 652 385 668
rect 232 603 234 607
rect 238 603 241 607
rect 245 603 248 607
rect 102 552 105 558
rect 182 552 185 558
rect 222 552 225 568
rect 94 542 97 548
rect 142 542 145 548
rect 82 538 86 541
rect 194 538 198 541
rect 122 528 126 531
rect 158 522 161 538
rect 46 472 49 488
rect 54 462 57 518
rect 78 471 81 518
rect 110 472 113 518
rect 166 512 169 518
rect 190 502 193 538
rect 198 502 201 528
rect 118 472 121 498
rect 126 482 129 488
rect 78 468 86 471
rect 26 458 30 461
rect 66 458 70 461
rect 6 442 9 448
rect 38 372 41 458
rect 66 448 70 451
rect 66 358 70 361
rect 78 352 81 358
rect 62 342 65 348
rect 86 342 89 468
rect 142 462 145 478
rect 150 462 153 468
rect 158 462 161 468
rect 166 462 169 488
rect 174 472 177 478
rect 106 458 110 461
rect 118 452 121 458
rect 94 432 97 448
rect 94 342 97 348
rect 6 272 9 338
rect 54 302 57 338
rect 86 332 89 338
rect 62 312 65 318
rect 54 292 57 298
rect 66 288 70 291
rect 54 272 57 288
rect 78 272 81 278
rect 66 248 70 251
rect 38 182 41 218
rect 38 162 41 168
rect 54 162 57 188
rect 62 152 65 178
rect 70 152 73 158
rect 50 148 54 151
rect 6 142 9 148
rect 66 138 70 141
rect 78 92 81 268
rect 86 252 89 308
rect 94 252 97 338
rect 102 262 105 428
rect 118 362 121 448
rect 182 382 185 478
rect 110 342 113 358
rect 118 352 121 358
rect 118 332 121 338
rect 110 241 113 318
rect 118 272 121 288
rect 106 238 113 241
rect 126 262 129 368
rect 162 348 166 351
rect 182 341 185 378
rect 178 338 185 341
rect 190 342 193 478
rect 198 452 201 498
rect 206 482 209 518
rect 230 482 233 538
rect 238 532 241 538
rect 246 522 249 548
rect 254 532 257 618
rect 342 592 345 618
rect 350 592 353 618
rect 230 472 233 478
rect 218 468 222 471
rect 206 462 209 468
rect 232 403 234 407
rect 238 403 241 407
rect 245 403 248 407
rect 254 392 257 468
rect 262 452 265 538
rect 270 532 273 558
rect 278 542 281 548
rect 270 372 273 528
rect 326 522 329 538
rect 294 482 297 518
rect 306 468 310 471
rect 286 462 289 468
rect 278 452 281 458
rect 302 452 305 458
rect 310 452 313 458
rect 318 452 321 458
rect 202 358 206 361
rect 242 358 246 361
rect 206 352 209 358
rect 142 322 145 328
rect 150 282 153 328
rect 146 278 150 281
rect 166 262 169 278
rect 182 262 185 288
rect 94 192 97 218
rect 94 132 97 168
rect 110 142 113 178
rect 126 152 129 258
rect 150 252 153 258
rect 134 182 137 238
rect 142 232 145 248
rect 134 152 137 178
rect 126 142 129 148
rect 30 72 33 78
rect 78 72 81 88
rect 94 71 97 128
rect 90 68 97 71
rect 134 70 137 98
rect 142 72 145 188
rect 150 162 153 218
rect 182 192 185 218
rect 162 148 166 151
rect 182 142 185 178
rect 190 172 193 338
rect 198 282 201 318
rect 206 312 209 338
rect 206 272 209 278
rect 198 252 201 258
rect 206 182 209 268
rect 214 262 217 348
rect 222 292 225 318
rect 230 262 233 328
rect 254 252 257 368
rect 286 352 289 358
rect 286 332 289 338
rect 302 332 305 418
rect 310 352 313 358
rect 326 352 329 518
rect 334 462 337 588
rect 358 542 361 568
rect 342 492 345 538
rect 366 512 369 548
rect 374 542 377 638
rect 390 542 393 548
rect 406 542 409 688
rect 462 672 465 678
rect 434 668 438 671
rect 414 652 417 658
rect 422 641 425 668
rect 442 658 446 661
rect 466 658 470 661
rect 454 652 457 658
rect 414 638 425 641
rect 438 642 441 648
rect 414 632 417 638
rect 406 532 409 538
rect 366 472 369 498
rect 354 468 358 471
rect 374 462 377 508
rect 398 472 401 488
rect 414 482 417 628
rect 422 531 425 578
rect 430 562 433 618
rect 438 562 441 588
rect 454 562 457 588
rect 474 548 478 551
rect 434 538 438 541
rect 422 528 433 531
rect 410 478 414 481
rect 422 472 425 518
rect 430 492 433 528
rect 454 472 457 518
rect 462 482 465 528
rect 470 512 473 518
rect 486 482 489 668
rect 494 662 497 678
rect 502 662 505 668
rect 502 532 505 558
rect 518 542 521 728
rect 534 728 538 732
rect 630 728 634 732
rect 710 728 714 732
rect 774 731 778 732
rect 774 728 785 731
rect 534 702 537 728
rect 608 703 610 707
rect 614 703 617 707
rect 621 703 624 707
rect 534 662 537 668
rect 550 662 553 678
rect 526 652 529 658
rect 558 602 561 618
rect 526 562 529 568
rect 538 558 542 561
rect 530 548 534 551
rect 566 542 569 698
rect 630 682 633 728
rect 710 702 713 728
rect 630 672 633 678
rect 670 672 673 678
rect 734 672 737 698
rect 782 692 785 728
rect 794 678 798 681
rect 586 668 590 671
rect 682 668 686 671
rect 734 662 737 668
rect 578 658 582 661
rect 594 658 598 661
rect 658 658 662 661
rect 750 652 753 658
rect 682 648 686 651
rect 586 568 590 571
rect 598 562 601 618
rect 606 562 609 568
rect 590 542 593 548
rect 514 538 518 541
rect 526 532 529 538
rect 494 492 497 518
rect 502 482 505 528
rect 522 478 526 481
rect 422 462 425 468
rect 454 462 457 468
rect 462 462 465 478
rect 526 462 529 468
rect 474 458 478 461
rect 498 458 502 461
rect 338 448 350 451
rect 374 351 377 458
rect 390 452 393 458
rect 418 428 422 431
rect 478 402 481 418
rect 370 348 377 351
rect 406 352 409 358
rect 262 322 265 328
rect 270 302 273 328
rect 286 282 289 298
rect 302 282 305 328
rect 318 292 321 318
rect 326 281 329 338
rect 342 332 345 338
rect 358 322 361 338
rect 318 278 329 281
rect 274 268 278 271
rect 286 262 289 278
rect 318 272 321 278
rect 314 268 318 271
rect 326 262 329 268
rect 334 262 337 288
rect 206 152 209 158
rect 178 128 182 131
rect 190 121 193 148
rect 198 132 201 138
rect 214 132 217 218
rect 232 203 234 207
rect 238 203 241 207
rect 245 203 248 207
rect 254 182 257 248
rect 222 162 225 168
rect 254 162 257 178
rect 230 152 233 158
rect 242 148 246 151
rect 182 118 193 121
rect 150 72 153 118
rect 166 102 169 118
rect 182 92 185 118
rect 238 92 241 108
rect 182 75 186 78
rect 254 72 257 78
rect 270 72 273 148
rect 278 82 281 138
rect 286 92 289 148
rect 294 142 297 218
rect 310 192 313 228
rect 334 222 337 258
rect 326 162 329 168
rect 342 162 345 318
rect 366 302 369 328
rect 350 282 353 288
rect 366 272 369 298
rect 374 272 377 348
rect 382 332 385 338
rect 406 332 409 338
rect 398 322 401 328
rect 382 272 385 318
rect 406 311 409 328
rect 398 308 409 311
rect 398 282 401 308
rect 358 262 361 268
rect 350 192 353 248
rect 366 162 369 218
rect 382 211 385 268
rect 390 262 393 268
rect 398 262 401 278
rect 374 208 385 211
rect 322 148 326 151
rect 310 132 313 138
rect 318 122 321 138
rect 358 132 361 138
rect 310 118 318 121
rect 310 92 313 118
rect 342 92 345 98
rect 302 72 305 78
rect 318 72 321 78
rect 366 72 369 128
rect 374 102 377 208
rect 386 158 390 161
rect 382 122 385 148
rect 390 142 393 148
rect 398 112 401 258
rect 414 242 417 258
rect 422 241 425 358
rect 430 342 433 378
rect 450 358 454 361
rect 486 342 489 348
rect 454 322 457 328
rect 470 322 473 338
rect 494 302 497 458
rect 534 452 537 518
rect 550 462 553 528
rect 558 472 561 538
rect 566 532 569 538
rect 574 482 577 538
rect 574 472 577 478
rect 562 468 566 471
rect 542 362 545 458
rect 582 452 585 528
rect 598 512 601 548
rect 614 522 617 638
rect 710 622 713 628
rect 742 622 745 648
rect 758 632 761 668
rect 806 652 809 658
rect 734 618 742 621
rect 646 562 649 568
rect 626 558 630 561
rect 622 522 625 528
rect 608 503 610 507
rect 614 503 617 507
rect 621 503 624 507
rect 598 462 601 468
rect 566 392 569 418
rect 598 392 601 418
rect 622 412 625 438
rect 558 372 561 378
rect 538 348 542 351
rect 554 348 558 351
rect 502 332 505 348
rect 566 342 569 378
rect 574 342 577 358
rect 602 348 606 351
rect 590 342 593 348
rect 502 312 505 328
rect 494 292 497 298
rect 446 282 449 288
rect 510 282 513 338
rect 518 332 521 338
rect 598 332 601 348
rect 622 342 625 408
rect 630 362 633 518
rect 638 492 641 548
rect 662 542 665 548
rect 670 542 673 598
rect 678 552 681 558
rect 698 548 702 551
rect 710 542 713 618
rect 734 592 737 618
rect 718 562 721 568
rect 690 538 694 541
rect 714 538 718 541
rect 650 528 654 531
rect 654 472 657 488
rect 702 472 705 518
rect 726 472 729 548
rect 734 522 737 548
rect 750 542 753 548
rect 758 542 761 618
rect 806 592 809 618
rect 822 582 825 618
rect 814 552 817 558
rect 822 552 825 568
rect 846 562 849 678
rect 870 582 873 588
rect 806 542 809 548
rect 778 538 782 541
rect 794 538 798 541
rect 742 522 745 538
rect 646 462 649 468
rect 674 458 678 461
rect 638 452 641 458
rect 662 362 665 458
rect 686 392 689 468
rect 694 382 697 418
rect 670 352 673 368
rect 694 352 697 378
rect 710 352 713 448
rect 718 412 721 458
rect 726 452 729 458
rect 718 362 721 408
rect 682 348 686 351
rect 538 328 542 331
rect 646 322 649 348
rect 586 318 590 321
rect 518 282 521 288
rect 506 278 510 281
rect 430 272 433 278
rect 562 268 566 271
rect 578 268 582 271
rect 454 252 457 268
rect 466 258 478 261
rect 482 258 486 261
rect 494 252 497 268
rect 546 258 550 261
rect 590 261 593 318
rect 598 282 601 308
rect 608 303 610 307
rect 614 303 617 307
rect 621 303 624 307
rect 634 278 638 281
rect 638 272 641 278
rect 654 272 657 348
rect 694 342 697 348
rect 682 338 686 341
rect 722 338 726 341
rect 670 332 673 338
rect 682 328 686 331
rect 734 291 737 488
rect 750 471 753 538
rect 822 532 825 538
rect 774 492 777 528
rect 782 522 785 528
rect 778 478 782 481
rect 750 468 761 471
rect 746 458 750 461
rect 758 452 761 468
rect 790 462 793 518
rect 814 492 817 528
rect 830 492 833 558
rect 846 532 849 548
rect 850 488 854 491
rect 822 482 825 488
rect 798 472 801 478
rect 866 468 870 471
rect 846 462 849 468
rect 774 442 777 448
rect 782 442 785 458
rect 814 452 817 458
rect 742 422 745 438
rect 750 432 753 438
rect 790 432 793 448
rect 758 372 761 418
rect 742 362 745 368
rect 774 362 777 428
rect 822 402 825 418
rect 802 368 806 371
rect 762 348 766 351
rect 742 342 745 348
rect 774 322 777 358
rect 790 342 793 348
rect 814 342 817 378
rect 822 362 825 368
rect 830 351 833 388
rect 838 362 841 398
rect 846 382 849 458
rect 854 452 857 468
rect 854 352 857 448
rect 830 348 841 351
rect 802 338 806 341
rect 730 288 737 291
rect 774 292 777 298
rect 738 278 742 281
rect 686 272 689 278
rect 646 262 649 268
rect 694 262 697 278
rect 730 268 734 271
rect 738 268 745 271
rect 762 268 766 271
rect 710 262 713 268
rect 582 258 593 261
rect 418 238 425 241
rect 478 242 481 248
rect 514 238 518 241
rect 446 202 449 218
rect 410 148 414 151
rect 446 142 449 158
rect 454 152 457 168
rect 462 162 465 218
rect 478 142 481 158
rect 498 148 502 151
rect 414 112 417 138
rect 438 132 441 140
rect 454 132 457 138
rect 474 128 478 131
rect 486 122 489 148
rect 510 142 513 218
rect 526 162 529 218
rect 558 192 561 218
rect 534 152 537 158
rect 494 132 497 138
rect 414 82 417 88
rect 422 72 425 118
rect 274 68 278 71
rect 206 62 209 68
rect 26 58 30 61
rect 106 58 110 61
rect 6 42 9 48
rect 232 3 234 7
rect 238 3 241 7
rect 245 3 248 7
rect 302 -18 305 68
rect 326 62 329 68
rect 326 -18 329 58
rect 374 52 377 68
rect 414 62 417 68
rect 438 62 441 88
rect 446 72 449 98
rect 458 78 462 81
rect 470 72 473 88
rect 510 82 513 108
rect 518 92 521 148
rect 542 142 545 178
rect 554 158 558 161
rect 566 152 569 258
rect 574 172 577 178
rect 582 152 585 258
rect 614 252 617 258
rect 530 138 534 141
rect 550 112 553 148
rect 590 142 593 248
rect 626 148 630 151
rect 638 142 641 258
rect 582 122 585 138
rect 526 92 529 108
rect 558 92 561 118
rect 590 112 593 138
rect 598 122 601 140
rect 646 122 649 258
rect 662 252 665 258
rect 670 242 673 248
rect 694 212 697 248
rect 608 103 610 107
rect 614 103 617 107
rect 621 103 624 107
rect 630 92 633 118
rect 630 82 633 88
rect 510 72 513 78
rect 542 72 545 78
rect 598 72 601 78
rect 606 72 609 78
rect 654 72 657 198
rect 662 152 665 158
rect 670 152 673 208
rect 686 152 689 158
rect 706 148 710 151
rect 718 142 721 188
rect 742 152 745 268
rect 790 152 793 278
rect 798 242 801 248
rect 806 202 809 268
rect 814 262 817 278
rect 822 272 825 348
rect 838 272 841 348
rect 846 342 849 348
rect 826 248 830 251
rect 838 202 841 268
rect 846 222 849 258
rect 862 252 865 418
rect 870 342 873 348
rect 830 162 833 168
rect 802 158 806 161
rect 846 152 849 218
rect 854 192 857 218
rect 862 152 865 198
rect 802 148 806 151
rect 826 148 830 151
rect 774 142 777 148
rect 674 138 678 141
rect 694 132 697 138
rect 750 132 753 138
rect 710 122 713 128
rect 666 118 670 121
rect 718 92 721 128
rect 766 122 769 128
rect 738 118 742 121
rect 758 112 761 118
rect 774 102 777 138
rect 450 68 457 71
rect 482 68 486 71
rect 610 68 614 71
rect 394 58 398 61
rect 422 52 425 58
rect 454 52 457 68
rect 526 62 529 68
rect 498 58 502 61
rect 542 52 545 68
rect 302 -22 306 -18
rect 326 -22 330 -18
rect 350 -19 353 18
rect 550 -18 553 38
rect 574 -18 577 68
rect 630 62 633 68
rect 662 62 665 78
rect 678 52 681 88
rect 734 72 737 98
rect 782 92 785 148
rect 862 142 865 148
rect 826 138 830 141
rect 790 72 793 98
rect 798 82 801 138
rect 842 128 846 131
rect 742 62 745 68
rect 814 62 817 68
rect 794 58 798 61
rect 838 52 841 108
rect 642 48 646 51
rect 674 48 678 51
rect 358 -19 362 -18
rect 350 -22 362 -19
rect 550 -22 554 -18
rect 574 -22 578 -18
rect 854 -19 858 -18
rect 862 -19 865 18
rect 854 -22 865 -19
<< m3contact >>
rect 38 698 42 702
rect 150 698 154 702
rect 326 698 330 702
rect 342 698 346 702
rect 302 688 306 692
rect 206 678 210 682
rect 238 678 242 682
rect 30 668 34 672
rect 6 648 10 652
rect 54 648 58 652
rect 14 558 18 562
rect 46 558 50 562
rect 6 548 10 552
rect 14 548 18 552
rect 30 548 34 552
rect 22 528 26 532
rect 6 518 10 522
rect 54 538 58 542
rect 94 668 98 672
rect 102 658 106 662
rect 126 658 130 662
rect 86 648 90 652
rect 110 628 114 632
rect 126 578 130 582
rect 78 568 82 572
rect 174 668 178 672
rect 166 648 170 652
rect 190 638 194 642
rect 318 678 322 682
rect 358 688 362 692
rect 406 688 410 692
rect 254 668 258 672
rect 334 668 338 672
rect 254 658 258 662
rect 310 658 314 662
rect 222 628 226 632
rect 294 648 298 652
rect 382 678 386 682
rect 390 668 394 672
rect 374 658 378 662
rect 310 638 314 642
rect 342 638 346 642
rect 374 638 378 642
rect 270 618 274 622
rect 342 618 346 622
rect 234 603 238 607
rect 241 603 245 607
rect 150 588 154 592
rect 222 568 226 572
rect 102 558 106 562
rect 142 558 146 562
rect 182 558 186 562
rect 78 538 82 542
rect 94 538 98 542
rect 142 538 146 542
rect 198 538 202 542
rect 230 538 234 542
rect 238 538 242 542
rect 62 528 66 532
rect 118 528 122 532
rect 158 518 162 522
rect 46 488 50 492
rect 166 508 170 512
rect 118 498 122 502
rect 190 498 194 502
rect 198 498 202 502
rect 166 488 170 492
rect 126 478 130 482
rect 142 478 146 482
rect 110 468 114 472
rect 30 458 34 462
rect 70 458 74 462
rect 6 448 10 452
rect 70 448 74 452
rect 38 368 42 372
rect 70 358 74 362
rect 78 358 82 362
rect 174 478 178 482
rect 182 478 186 482
rect 102 458 106 462
rect 118 458 122 462
rect 150 458 154 462
rect 158 458 162 462
rect 166 458 170 462
rect 118 448 122 452
rect 94 428 98 432
rect 102 428 106 432
rect 94 348 98 352
rect 62 338 66 342
rect 86 328 90 332
rect 62 308 66 312
rect 86 308 90 312
rect 54 298 58 302
rect 54 288 58 292
rect 62 288 66 292
rect 78 278 82 282
rect 6 268 10 272
rect 70 248 74 252
rect 54 188 58 192
rect 38 178 42 182
rect 62 178 66 182
rect 38 158 42 162
rect 6 148 10 152
rect 54 148 58 152
rect 70 148 74 152
rect 70 138 74 142
rect 182 378 186 382
rect 126 368 130 372
rect 118 358 122 362
rect 110 338 114 342
rect 118 328 122 332
rect 102 258 106 262
rect 94 248 98 252
rect 118 288 122 292
rect 158 348 162 352
rect 174 338 178 342
rect 238 528 242 532
rect 334 588 338 592
rect 350 588 354 592
rect 254 528 258 532
rect 246 518 250 522
rect 206 478 210 482
rect 230 478 234 482
rect 222 468 226 472
rect 206 458 210 462
rect 198 448 202 452
rect 234 403 238 407
rect 241 403 245 407
rect 278 548 282 552
rect 270 528 274 532
rect 262 448 266 452
rect 254 388 258 392
rect 326 518 330 522
rect 294 478 298 482
rect 286 468 290 472
rect 302 468 306 472
rect 278 458 282 462
rect 318 458 322 462
rect 302 448 306 452
rect 310 448 314 452
rect 302 418 306 422
rect 254 368 258 372
rect 270 368 274 372
rect 206 358 210 362
rect 238 358 242 362
rect 214 348 218 352
rect 190 338 194 342
rect 142 328 146 332
rect 182 288 186 292
rect 142 278 146 282
rect 166 278 170 282
rect 94 188 98 192
rect 110 178 114 182
rect 94 168 98 172
rect 150 248 154 252
rect 134 238 138 242
rect 142 228 146 232
rect 150 218 154 222
rect 142 188 146 192
rect 134 178 138 182
rect 126 138 130 142
rect 78 88 82 92
rect 30 78 34 82
rect 134 98 138 102
rect 182 188 186 192
rect 182 178 186 182
rect 166 148 170 152
rect 206 308 210 312
rect 198 278 202 282
rect 206 278 210 282
rect 198 258 202 262
rect 222 288 226 292
rect 230 258 234 262
rect 286 358 290 362
rect 358 568 362 572
rect 390 548 394 552
rect 462 678 466 682
rect 494 678 498 682
rect 438 668 442 672
rect 486 668 490 672
rect 414 658 418 662
rect 446 658 450 662
rect 462 658 466 662
rect 454 648 458 652
rect 438 638 442 642
rect 414 628 418 632
rect 406 538 410 542
rect 366 508 370 512
rect 374 508 378 512
rect 366 498 370 502
rect 342 488 346 492
rect 358 468 362 472
rect 398 488 402 492
rect 422 578 426 582
rect 438 588 442 592
rect 454 588 458 592
rect 430 558 434 562
rect 470 548 474 552
rect 430 538 434 542
rect 414 478 418 482
rect 470 508 474 512
rect 502 658 506 662
rect 502 558 506 562
rect 610 703 614 707
rect 617 703 621 707
rect 534 698 538 702
rect 566 698 570 702
rect 534 668 538 672
rect 526 648 530 652
rect 558 598 562 602
rect 526 558 530 562
rect 534 558 538 562
rect 534 548 538 552
rect 710 698 714 702
rect 734 698 738 702
rect 670 678 674 682
rect 798 678 802 682
rect 846 678 850 682
rect 582 668 586 672
rect 630 668 634 672
rect 678 668 682 672
rect 582 658 586 662
rect 598 658 602 662
rect 654 658 658 662
rect 734 658 738 662
rect 750 658 754 662
rect 686 648 690 652
rect 590 568 594 572
rect 606 568 610 572
rect 598 558 602 562
rect 590 548 594 552
rect 598 548 602 552
rect 518 538 522 542
rect 558 538 562 542
rect 574 538 578 542
rect 526 528 530 532
rect 550 528 554 532
rect 494 488 498 492
rect 534 518 538 522
rect 462 478 466 482
rect 526 478 530 482
rect 422 468 426 472
rect 526 468 530 472
rect 390 458 394 462
rect 454 458 458 462
rect 470 458 474 462
rect 502 458 506 462
rect 310 348 314 352
rect 422 428 426 432
rect 478 398 482 402
rect 430 378 434 382
rect 406 358 410 362
rect 286 328 290 332
rect 262 318 266 322
rect 270 298 274 302
rect 286 298 290 302
rect 318 288 322 292
rect 342 328 346 332
rect 366 328 370 332
rect 358 318 362 322
rect 334 288 338 292
rect 270 268 274 272
rect 310 268 314 272
rect 326 258 330 262
rect 206 178 210 182
rect 190 168 194 172
rect 206 148 210 152
rect 182 128 186 132
rect 234 203 238 207
rect 241 203 245 207
rect 310 228 314 232
rect 254 178 258 182
rect 222 168 226 172
rect 230 158 234 162
rect 238 148 242 152
rect 198 128 202 132
rect 166 98 170 102
rect 238 108 242 112
rect 182 88 186 92
rect 182 78 186 82
rect 254 78 258 82
rect 334 218 338 222
rect 326 168 330 172
rect 366 298 370 302
rect 350 278 354 282
rect 382 328 386 332
rect 406 328 410 332
rect 382 318 386 322
rect 398 318 402 322
rect 358 268 362 272
rect 374 268 378 272
rect 390 268 394 272
rect 398 258 402 262
rect 366 158 370 162
rect 318 148 322 152
rect 310 138 314 142
rect 358 138 362 142
rect 318 118 322 122
rect 342 98 346 102
rect 278 78 282 82
rect 302 78 306 82
rect 318 78 322 82
rect 382 158 386 162
rect 390 138 394 142
rect 382 118 386 122
rect 414 238 418 242
rect 446 358 450 362
rect 486 348 490 352
rect 454 318 458 322
rect 470 318 474 322
rect 566 528 570 532
rect 582 528 586 532
rect 574 478 578 482
rect 566 468 570 472
rect 710 628 714 632
rect 806 648 810 652
rect 758 628 762 632
rect 742 618 746 622
rect 758 618 762 622
rect 670 598 674 602
rect 622 558 626 562
rect 646 558 650 562
rect 662 548 666 552
rect 614 518 618 522
rect 622 518 626 522
rect 630 518 634 522
rect 598 508 602 512
rect 610 503 614 507
rect 617 503 621 507
rect 598 468 602 472
rect 598 418 602 422
rect 622 408 626 412
rect 566 388 570 392
rect 558 378 562 382
rect 566 378 570 382
rect 534 348 538 352
rect 550 348 554 352
rect 574 358 578 362
rect 590 348 594 352
rect 606 348 610 352
rect 510 338 514 342
rect 502 308 506 312
rect 494 298 498 302
rect 446 288 450 292
rect 494 288 498 292
rect 678 558 682 562
rect 694 548 698 552
rect 718 568 722 572
rect 726 548 730 552
rect 686 538 690 542
rect 718 538 722 542
rect 646 528 650 532
rect 702 518 706 522
rect 654 488 658 492
rect 806 588 810 592
rect 822 578 826 582
rect 822 568 826 572
rect 814 558 818 562
rect 870 578 874 582
rect 846 558 850 562
rect 750 538 754 542
rect 782 538 786 542
rect 790 538 794 542
rect 806 538 810 542
rect 822 538 826 542
rect 734 518 738 522
rect 742 518 746 522
rect 734 488 738 492
rect 646 468 650 472
rect 638 458 642 462
rect 670 458 674 462
rect 718 458 722 462
rect 686 388 690 392
rect 694 378 698 382
rect 670 368 674 372
rect 726 448 730 452
rect 718 408 722 412
rect 654 348 658 352
rect 678 348 682 352
rect 518 328 522 332
rect 542 328 546 332
rect 598 328 602 332
rect 590 318 594 322
rect 646 318 650 322
rect 518 288 522 292
rect 430 278 434 282
rect 502 278 506 282
rect 558 268 562 272
rect 582 268 586 272
rect 478 258 482 262
rect 550 258 554 262
rect 598 308 602 312
rect 610 303 614 307
rect 617 303 621 307
rect 638 278 642 282
rect 678 338 682 342
rect 694 338 698 342
rect 718 338 722 342
rect 670 328 674 332
rect 678 328 682 332
rect 726 288 730 292
rect 814 528 818 532
rect 782 518 786 522
rect 774 488 778 492
rect 782 478 786 482
rect 742 458 746 462
rect 846 528 850 532
rect 822 488 826 492
rect 830 488 834 492
rect 846 488 850 492
rect 798 478 802 482
rect 846 468 850 472
rect 862 468 866 472
rect 790 458 794 462
rect 814 458 818 462
rect 774 448 778 452
rect 750 438 754 442
rect 782 438 786 442
rect 774 428 778 432
rect 790 428 794 432
rect 742 418 746 422
rect 758 418 762 422
rect 742 368 746 372
rect 822 398 826 402
rect 838 398 842 402
rect 830 388 834 392
rect 814 378 818 382
rect 806 368 810 372
rect 742 348 746 352
rect 758 348 762 352
rect 822 358 826 362
rect 822 348 826 352
rect 846 378 850 382
rect 862 418 866 422
rect 790 338 794 342
rect 798 338 802 342
rect 774 318 778 322
rect 774 298 778 302
rect 686 278 690 282
rect 694 278 698 282
rect 734 278 738 282
rect 814 278 818 282
rect 646 268 650 272
rect 726 268 730 272
rect 758 268 762 272
rect 638 258 642 262
rect 662 258 666 262
rect 710 258 714 262
rect 454 248 458 252
rect 494 248 498 252
rect 478 238 482 242
rect 510 238 514 242
rect 510 218 514 222
rect 446 198 450 202
rect 454 168 458 172
rect 446 158 450 162
rect 414 148 418 152
rect 462 158 466 162
rect 478 158 482 162
rect 494 148 498 152
rect 454 138 458 142
rect 438 128 442 132
rect 478 128 482 132
rect 558 188 562 192
rect 542 178 546 182
rect 526 158 530 162
rect 534 158 538 162
rect 494 128 498 132
rect 486 118 490 122
rect 398 108 402 112
rect 414 108 418 112
rect 374 98 378 102
rect 414 88 418 92
rect 510 108 514 112
rect 446 98 450 102
rect 438 88 442 92
rect 150 68 154 72
rect 206 68 210 72
rect 270 68 274 72
rect 326 68 330 72
rect 366 68 370 72
rect 374 68 378 72
rect 422 68 426 72
rect 30 58 34 62
rect 102 58 106 62
rect 6 48 10 52
rect 234 3 238 7
rect 241 3 245 7
rect 470 88 474 92
rect 462 78 466 82
rect 550 158 554 162
rect 574 178 578 182
rect 614 248 618 252
rect 566 148 570 152
rect 582 148 586 152
rect 534 138 538 142
rect 542 138 546 142
rect 622 148 626 152
rect 558 118 562 122
rect 582 118 586 122
rect 526 108 530 112
rect 550 108 554 112
rect 670 238 674 242
rect 670 208 674 212
rect 694 208 698 212
rect 654 198 658 202
rect 598 118 602 122
rect 646 118 650 122
rect 590 108 594 112
rect 610 103 614 107
rect 617 103 621 107
rect 518 88 522 92
rect 630 88 634 92
rect 510 78 514 82
rect 606 78 610 82
rect 630 78 634 82
rect 718 188 722 192
rect 686 158 690 162
rect 662 148 666 152
rect 710 148 714 152
rect 798 238 802 242
rect 854 348 858 352
rect 846 338 850 342
rect 822 248 826 252
rect 846 258 850 262
rect 870 348 874 352
rect 854 218 858 222
rect 806 198 810 202
rect 838 198 842 202
rect 806 158 810 162
rect 830 158 834 162
rect 862 198 866 202
rect 774 148 778 152
rect 806 148 810 152
rect 830 148 834 152
rect 846 148 850 152
rect 862 148 866 152
rect 670 138 674 142
rect 694 128 698 132
rect 718 128 722 132
rect 750 128 754 132
rect 670 118 674 122
rect 710 118 714 122
rect 742 118 746 122
rect 766 118 770 122
rect 758 108 762 112
rect 734 98 738 102
rect 774 98 778 102
rect 678 88 682 92
rect 662 78 666 82
rect 478 68 482 72
rect 542 68 546 72
rect 598 68 602 72
rect 614 68 618 72
rect 630 68 634 72
rect 398 58 402 62
rect 414 58 418 62
rect 422 58 426 62
rect 502 58 506 62
rect 526 58 530 62
rect 798 138 802 142
rect 822 138 826 142
rect 790 98 794 102
rect 782 88 786 92
rect 838 128 842 132
rect 838 108 842 112
rect 742 58 746 62
rect 798 58 802 62
rect 814 58 818 62
rect 646 48 650 52
rect 670 48 674 52
<< metal3 >>
rect 608 703 610 707
rect 614 703 617 707
rect 622 703 624 707
rect 42 698 150 701
rect 330 698 342 701
rect 538 698 566 701
rect 714 698 734 701
rect 306 688 358 691
rect 362 688 406 691
rect 210 678 238 681
rect 242 678 318 681
rect 322 678 382 681
rect 466 678 494 681
rect 498 678 670 681
rect 802 678 846 681
rect 34 668 94 671
rect 178 668 254 671
rect 338 668 377 671
rect 394 668 438 671
rect 490 668 505 671
rect 374 662 377 668
rect 502 662 505 668
rect 586 668 630 671
rect 634 668 646 671
rect 650 668 678 671
rect 106 658 126 661
rect 258 658 310 661
rect 450 658 462 661
rect 534 661 537 668
rect 506 658 537 661
rect 586 658 598 661
rect 602 658 654 661
rect 658 658 734 661
rect -26 651 -22 652
rect -26 648 6 651
rect 10 648 54 651
rect 58 648 86 651
rect 90 648 166 651
rect 414 651 417 658
rect 298 648 409 651
rect 414 648 454 651
rect 530 648 542 651
rect 750 651 753 658
rect 690 648 753 651
rect 806 652 809 658
rect 110 638 190 641
rect 314 638 342 641
rect 346 638 374 641
rect 406 641 409 648
rect 406 638 438 641
rect 110 632 113 638
rect 226 628 414 631
rect 714 628 758 631
rect 274 618 342 621
rect 746 618 758 621
rect 232 603 234 607
rect 238 603 241 607
rect 246 603 248 607
rect 562 598 670 601
rect 154 588 334 591
rect 354 588 438 591
rect 442 588 454 591
rect 810 588 846 591
rect 130 578 422 581
rect 826 578 830 581
rect 902 581 906 582
rect 874 578 906 581
rect 82 568 110 571
rect 114 568 222 571
rect 226 568 358 571
rect 594 568 606 571
rect 610 568 718 571
rect 722 568 822 571
rect 18 558 46 561
rect 146 558 182 561
rect 434 558 502 561
rect 530 558 534 561
rect 602 558 622 561
rect 650 558 678 561
rect 850 558 870 561
rect 902 561 906 562
rect 874 558 906 561
rect -26 551 -22 552
rect -26 548 6 551
rect 18 548 30 551
rect 102 551 105 558
rect 34 548 105 551
rect 394 548 470 551
rect 538 548 590 551
rect 602 548 662 551
rect 698 548 726 551
rect 814 551 817 558
rect 730 548 817 551
rect 58 538 78 541
rect 98 538 142 541
rect 202 538 230 541
rect 278 541 281 548
rect 242 538 281 541
rect 410 538 430 541
rect 522 538 558 541
rect 578 538 686 541
rect 722 538 750 541
rect 786 538 790 541
rect 810 538 822 541
rect -26 531 -22 532
rect -26 528 22 531
rect 26 528 62 531
rect 66 528 118 531
rect 122 528 238 531
rect 258 528 270 531
rect 274 528 345 531
rect 530 528 550 531
rect 554 528 566 531
rect 570 528 582 531
rect 650 528 785 531
rect 818 528 846 531
rect 10 518 158 521
rect 162 518 246 521
rect 250 518 326 521
rect 342 521 345 528
rect 782 522 785 528
rect 342 518 534 521
rect 538 518 614 521
rect 626 518 630 521
rect 634 518 702 521
rect 706 518 734 521
rect 746 518 750 521
rect 170 508 358 511
rect 370 508 374 511
rect 378 508 470 511
rect 474 508 574 511
rect 578 508 598 511
rect 608 503 610 507
rect 614 503 617 507
rect 622 503 624 507
rect 122 498 190 501
rect 202 498 366 501
rect 50 488 166 491
rect 346 488 398 491
rect 402 488 494 491
rect 498 488 654 491
rect 738 488 774 491
rect 778 488 822 491
rect 834 488 846 491
rect 66 478 126 481
rect 146 478 174 481
rect 186 478 206 481
rect 234 478 294 481
rect 418 478 462 481
rect 530 478 574 481
rect 786 478 798 481
rect 646 472 649 478
rect 114 468 121 471
rect 118 462 121 468
rect 158 468 222 471
rect 242 468 286 471
rect 306 468 310 471
rect 354 468 358 471
rect 426 468 526 471
rect 570 468 598 471
rect 850 468 862 471
rect 150 462 153 468
rect 158 462 161 468
rect 34 458 70 461
rect 106 458 110 461
rect 170 458 206 461
rect 302 458 318 461
rect 458 458 470 461
rect 506 458 638 461
rect 642 458 670 461
rect 722 458 742 461
rect 794 458 814 461
rect -26 451 -22 452
rect -26 448 6 451
rect 66 448 70 451
rect 122 448 198 451
rect 278 451 281 458
rect 266 448 281 451
rect 302 452 305 458
rect 314 448 326 451
rect 390 451 393 458
rect 330 448 393 451
rect 546 448 726 451
rect 730 448 774 451
rect 754 438 782 441
rect 98 428 102 431
rect 106 428 422 431
rect 426 428 774 431
rect 778 428 790 431
rect 306 418 310 421
rect 602 418 742 421
rect 746 418 758 421
rect 866 418 870 421
rect 626 408 718 411
rect 232 403 234 407
rect 238 403 241 407
rect 246 403 248 407
rect 482 398 678 401
rect 826 398 838 401
rect 218 388 254 391
rect 258 388 558 391
rect 562 388 566 391
rect 690 388 830 391
rect 186 378 430 381
rect 570 378 694 381
rect 698 378 814 381
rect 818 378 846 381
rect 42 368 126 371
rect 258 368 270 371
rect 558 371 561 378
rect 558 368 670 371
rect 810 368 825 371
rect 66 358 70 361
rect 82 358 118 361
rect 210 358 238 361
rect 290 358 313 361
rect 410 358 446 361
rect 578 358 582 361
rect 742 361 745 368
rect 690 358 745 361
rect 822 362 825 368
rect 310 352 313 358
rect 98 348 158 351
rect 162 348 214 351
rect 490 348 510 351
rect 538 348 542 351
rect 554 348 558 351
rect 586 348 590 351
rect 610 348 654 351
rect 682 348 737 351
rect 746 348 758 351
rect 826 348 854 351
rect 902 351 906 352
rect 874 348 906 351
rect 94 341 97 348
rect 66 338 97 341
rect 114 338 174 341
rect 194 338 510 341
rect 586 338 678 341
rect 682 338 686 341
rect 698 338 718 341
rect 734 341 737 348
rect 734 338 790 341
rect 802 338 846 341
rect 90 328 118 331
rect 262 328 286 331
rect 346 328 350 331
rect 354 328 366 331
rect 386 328 406 331
rect 454 328 518 331
rect 546 328 598 331
rect 674 328 678 331
rect 142 321 145 328
rect 262 322 265 328
rect 454 322 457 328
rect 142 318 246 321
rect 266 318 358 321
rect 386 318 398 321
rect 450 318 454 321
rect 466 318 470 321
rect 582 318 590 321
rect 594 318 646 321
rect 774 312 777 318
rect 66 308 86 311
rect 90 308 206 311
rect 506 308 598 311
rect 608 303 610 307
rect 614 303 617 307
rect 622 303 624 307
rect 58 298 270 301
rect 274 298 286 301
rect 370 298 494 301
rect 746 298 774 301
rect -26 291 -22 292
rect -26 288 54 291
rect 66 288 118 291
rect 186 288 222 291
rect 322 288 334 291
rect 350 288 446 291
rect 498 288 518 291
rect 526 288 726 291
rect 350 282 353 288
rect 82 278 142 281
rect 170 278 198 281
rect 210 278 214 281
rect 362 278 430 281
rect 526 281 529 288
rect 506 278 529 281
rect 642 278 686 281
rect 698 278 734 281
rect 738 278 814 281
rect -26 271 -22 272
rect -26 268 6 271
rect 10 268 270 271
rect 274 268 310 271
rect 314 268 358 271
rect 378 268 390 271
rect 538 268 558 271
rect 586 268 646 271
rect 682 268 726 271
rect 762 268 766 271
rect 106 258 198 261
rect 234 258 326 261
rect 330 258 398 261
rect 482 258 505 261
rect 546 258 550 261
rect 642 258 662 261
rect 666 258 710 261
rect 714 258 846 261
rect 74 248 94 251
rect 154 248 454 251
rect 458 248 494 251
rect 502 251 505 258
rect 502 248 614 251
rect 618 248 673 251
rect 670 242 673 248
rect 798 248 822 251
rect 798 242 801 248
rect 138 238 414 241
rect 482 238 510 241
rect 146 228 310 231
rect 154 218 334 221
rect 514 218 806 221
rect 810 218 854 221
rect 674 208 694 211
rect 698 208 830 211
rect 232 203 234 207
rect 238 203 241 207
rect 246 203 248 207
rect 450 198 654 201
rect 658 198 806 201
rect 842 198 862 201
rect 58 188 94 191
rect 146 188 182 191
rect 562 188 718 191
rect 42 178 62 181
rect 66 178 110 181
rect 114 178 134 181
rect 186 178 206 181
rect 258 178 542 181
rect 98 168 190 171
rect 574 171 577 178
rect 458 168 577 171
rect 222 161 225 168
rect 42 158 225 161
rect 326 161 329 168
rect 234 158 329 161
rect 370 158 382 161
rect 450 158 462 161
rect 482 158 526 161
rect 538 158 550 161
rect 662 158 686 161
rect 810 158 830 161
rect 662 152 665 158
rect -26 151 -22 152
rect -26 148 6 151
rect 58 148 70 151
rect 162 148 166 151
rect 210 148 238 151
rect 322 148 326 151
rect 330 148 414 151
rect 418 148 494 151
rect 498 148 566 151
rect 586 148 622 151
rect 714 148 774 151
rect 778 148 806 151
rect 834 148 846 151
rect 902 151 906 152
rect 866 148 906 151
rect 74 138 126 141
rect 370 138 390 141
rect 438 138 454 141
rect 530 138 534 141
rect 546 138 670 141
rect 778 138 798 141
rect 826 138 830 141
rect 186 128 198 131
rect 310 131 313 138
rect 358 131 361 138
rect 310 128 361 131
rect 438 132 441 138
rect 482 128 494 131
rect 534 131 537 138
rect 534 128 694 131
rect 722 128 750 131
rect 842 128 846 131
rect 322 118 382 121
rect 386 118 486 121
rect 562 118 582 121
rect 586 118 598 121
rect 602 118 646 121
rect 662 118 670 121
rect 674 118 710 121
rect 734 118 742 121
rect 746 118 766 121
rect 242 108 398 111
rect 418 108 510 111
rect 530 108 550 111
rect 554 108 590 111
rect 762 108 838 111
rect 608 103 610 107
rect 614 103 617 107
rect 622 103 624 107
rect 138 98 166 101
rect 346 98 374 101
rect 450 98 454 101
rect 738 98 774 101
rect 778 98 790 101
rect 82 88 182 91
rect 442 88 470 91
rect 474 88 518 91
rect 522 88 630 91
rect 682 88 782 91
rect 186 78 254 81
rect 258 78 278 81
rect 282 78 302 81
rect 306 78 318 81
rect 414 81 417 88
rect 414 78 462 81
rect 514 78 542 81
rect 546 78 606 81
rect 634 78 662 81
rect 30 71 33 78
rect 30 68 150 71
rect 210 68 270 71
rect 274 68 326 71
rect 330 68 366 71
rect 378 68 422 71
rect 482 68 537 71
rect 546 68 598 71
rect 618 68 630 71
rect 34 58 102 61
rect 402 58 414 61
rect 506 58 526 61
rect 534 61 537 68
rect 534 58 742 61
rect 802 58 814 61
rect 422 52 425 58
rect -26 51 -22 52
rect -26 48 6 51
rect 650 48 670 51
rect 232 3 234 7
rect 238 3 241 7
rect 246 3 248 7
<< m4contact >>
rect 610 703 614 707
rect 618 703 621 707
rect 621 703 622 707
rect 646 668 650 672
rect 806 658 810 662
rect 542 648 546 652
rect 234 603 238 607
rect 242 603 245 607
rect 245 603 246 607
rect 846 588 850 592
rect 830 578 834 582
rect 110 568 114 572
rect 534 558 538 562
rect 870 558 874 562
rect 750 518 754 522
rect 358 508 362 512
rect 574 508 578 512
rect 610 503 614 507
rect 618 503 621 507
rect 621 503 622 507
rect 62 478 66 482
rect 526 478 530 482
rect 646 478 650 482
rect 150 468 154 472
rect 238 468 242 472
rect 310 468 314 472
rect 350 468 354 472
rect 110 458 114 462
rect 62 448 66 452
rect 326 448 330 452
rect 542 448 546 452
rect 422 428 426 432
rect 310 418 314 422
rect 870 418 874 422
rect 234 403 238 407
rect 242 403 245 407
rect 245 403 246 407
rect 678 398 682 402
rect 214 388 218 392
rect 558 388 562 392
rect 62 358 66 362
rect 582 358 586 362
rect 686 358 690 362
rect 510 348 514 352
rect 542 348 546 352
rect 558 348 562 352
rect 582 348 586 352
rect 582 338 586 342
rect 686 338 690 342
rect 350 328 354 332
rect 246 318 250 322
rect 446 318 450 322
rect 462 318 466 322
rect 774 308 778 312
rect 610 303 614 307
rect 618 303 621 307
rect 621 303 622 307
rect 742 298 746 302
rect 214 278 218 282
rect 358 278 362 282
rect 534 268 538 272
rect 678 268 682 272
rect 766 268 770 272
rect 542 258 546 262
rect 494 248 498 252
rect 806 218 810 222
rect 830 208 834 212
rect 234 203 238 207
rect 242 203 245 207
rect 245 203 246 207
rect 62 178 66 182
rect 158 148 162 152
rect 326 148 330 152
rect 366 138 370 142
rect 526 138 530 142
rect 774 138 778 142
rect 830 138 834 142
rect 846 128 850 132
rect 610 103 614 107
rect 618 103 621 107
rect 621 103 622 107
rect 454 98 458 102
rect 542 78 546 82
rect 422 48 426 52
rect 234 3 238 7
rect 242 3 245 7
rect 245 3 246 7
<< metal4 >>
rect 608 703 610 707
rect 614 703 617 707
rect 622 703 624 707
rect 232 603 234 607
rect 238 603 241 607
rect 246 603 248 607
rect 62 452 65 478
rect 110 462 113 568
rect 154 468 158 471
rect 234 468 238 471
rect 310 422 313 468
rect 232 403 234 407
rect 238 403 241 407
rect 246 403 248 407
rect 62 182 65 358
rect 214 282 217 388
rect 250 318 254 321
rect 232 203 234 207
rect 238 203 241 207
rect 246 203 248 207
rect 326 152 329 448
rect 350 332 353 468
rect 358 282 361 508
rect 162 148 166 151
rect 366 142 369 148
rect 422 52 425 428
rect 514 348 518 351
rect 466 318 470 321
rect 446 101 449 318
rect 494 252 497 268
rect 526 142 529 478
rect 534 272 537 558
rect 542 452 545 648
rect 558 352 561 388
rect 574 361 577 508
rect 608 503 610 507
rect 614 503 617 507
rect 622 503 624 507
rect 646 482 649 668
rect 742 518 750 521
rect 574 358 582 361
rect 586 348 590 351
rect 542 342 545 348
rect 578 338 582 341
rect 608 303 610 307
rect 614 303 617 307
rect 622 303 624 307
rect 678 272 681 398
rect 686 342 689 358
rect 742 302 745 518
rect 762 268 766 271
rect 446 98 454 101
rect 542 82 545 258
rect 774 142 777 308
rect 806 222 809 658
rect 830 212 833 578
rect 830 142 833 208
rect 846 132 849 588
rect 870 422 873 558
rect 608 103 610 107
rect 614 103 617 107
rect 622 103 624 107
rect 232 3 234 7
rect 238 3 241 7
rect 246 3 248 7
<< m5contact >>
rect 610 703 614 707
rect 617 703 618 707
rect 618 703 621 707
rect 234 603 238 607
rect 241 603 242 607
rect 242 603 245 607
rect 158 468 162 472
rect 230 468 234 472
rect 234 403 238 407
rect 241 403 242 407
rect 242 403 245 407
rect 254 318 258 322
rect 234 203 238 207
rect 241 203 242 207
rect 242 203 245 207
rect 166 148 170 152
rect 366 148 370 152
rect 518 348 522 352
rect 470 318 474 322
rect 494 268 498 272
rect 610 503 614 507
rect 617 503 618 507
rect 618 503 621 507
rect 590 348 594 352
rect 542 338 546 342
rect 574 338 578 342
rect 610 303 614 307
rect 617 303 618 307
rect 618 303 621 307
rect 758 268 762 272
rect 610 103 614 107
rect 617 103 618 107
rect 618 103 621 107
rect 234 3 238 7
rect 241 3 242 7
rect 242 3 245 7
<< metal5 >>
rect 614 703 617 707
rect 613 702 618 703
rect 623 702 624 707
rect 238 603 241 607
rect 237 602 242 603
rect 247 602 248 607
rect 614 503 617 507
rect 613 502 618 503
rect 623 502 624 507
rect 162 468 230 471
rect 238 403 241 407
rect 237 402 242 403
rect 247 402 248 407
rect 522 348 590 351
rect 546 338 574 341
rect 258 318 470 321
rect 614 303 617 307
rect 613 302 618 303
rect 623 302 624 307
rect 498 268 758 271
rect 238 203 241 207
rect 237 202 242 203
rect 247 202 248 207
rect 170 148 366 151
rect 614 103 617 107
rect 613 102 618 103
rect 623 102 624 107
rect 238 3 241 7
rect 237 2 242 3
rect 247 2 248 7
<< m6contact >>
rect 608 703 610 707
rect 610 703 613 707
rect 618 703 621 707
rect 621 703 623 707
rect 608 702 613 703
rect 618 702 623 703
rect 232 603 234 607
rect 234 603 237 607
rect 242 603 245 607
rect 245 603 247 607
rect 232 602 237 603
rect 242 602 247 603
rect 608 503 610 507
rect 610 503 613 507
rect 618 503 621 507
rect 621 503 623 507
rect 608 502 613 503
rect 618 502 623 503
rect 232 403 234 407
rect 234 403 237 407
rect 242 403 245 407
rect 245 403 247 407
rect 232 402 237 403
rect 242 402 247 403
rect 608 303 610 307
rect 610 303 613 307
rect 618 303 621 307
rect 621 303 623 307
rect 608 302 613 303
rect 618 302 623 303
rect 232 203 234 207
rect 234 203 237 207
rect 242 203 245 207
rect 245 203 247 207
rect 232 202 237 203
rect 242 202 247 203
rect 608 103 610 107
rect 610 103 613 107
rect 618 103 621 107
rect 621 103 623 107
rect 608 102 613 103
rect 618 102 623 103
rect 232 3 234 7
rect 234 3 237 7
rect 242 3 245 7
rect 245 3 247 7
rect 232 2 237 3
rect 242 2 247 3
<< metal6 >>
rect 232 607 248 730
rect 237 602 242 607
rect 247 602 248 607
rect 232 407 248 602
rect 237 402 242 407
rect 247 402 248 407
rect 232 207 248 402
rect 237 202 242 207
rect 247 202 248 207
rect 232 7 248 202
rect 237 2 242 7
rect 247 2 248 7
rect 232 -30 248 2
rect 608 707 624 730
rect 613 702 618 707
rect 623 702 624 707
rect 608 507 624 702
rect 613 502 618 507
rect 623 502 624 507
rect 608 307 624 502
rect 613 302 618 307
rect 623 302 624 307
rect 608 107 624 302
rect 613 102 618 107
rect 623 102 624 107
rect 608 -30 624 102
use BUFX2  BUFX2_4
timestamp 1743078376
transform -1 0 28 0 -1 105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_4
timestamp 1743078376
transform 1 0 28 0 -1 105
box -2 -3 58 103
use BUFX2  BUFX2_3
timestamp 1743078376
transform -1 0 28 0 1 105
box -2 -3 26 103
use NAND3X1  NAND3X1_4
timestamp 1743078376
transform -1 0 60 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_22
timestamp 1743078376
transform 1 0 60 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_32
timestamp 1743078376
transform 1 0 84 0 -1 105
box -2 -3 34 103
use AND2X2  AND2X2_6
timestamp 1743078376
transform -1 0 148 0 -1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_11
timestamp 1743078376
transform -1 0 124 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_26
timestamp 1743078376
transform 1 0 124 0 1 105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_2
timestamp 1743078376
transform 1 0 148 0 -1 105
box -2 -3 58 103
use NOR2X1  NOR2X1_22
timestamp 1743078376
transform -1 0 180 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_30
timestamp 1743078376
transform 1 0 180 0 1 105
box -2 -3 34 103
use XOR2X1  XOR2X1_2
timestamp 1743078376
transform -1 0 260 0 -1 105
box -2 -3 58 103
use NOR2X1  NOR2X1_20
timestamp 1743078376
transform 1 0 212 0 1 105
box -2 -3 26 103
use FILL  FILL_1_0_0
timestamp 1743078376
transform -1 0 244 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_1
timestamp 1743078376
transform -1 0 252 0 1 105
box -2 -3 10 103
use FILL  FILL_0_0_0
timestamp 1743078376
transform 1 0 260 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1743078376
transform 1 0 268 0 -1 105
box -2 -3 10 103
use NAND2X1  NAND2X1_11
timestamp 1743078376
transform 1 0 276 0 -1 105
box -2 -3 26 103
use INVX2  INVX2_6
timestamp 1743078376
transform 1 0 300 0 -1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_29
timestamp 1743078376
transform -1 0 284 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_4
timestamp 1743078376
transform 1 0 284 0 1 105
box -2 -3 34 103
use AND2X2  AND2X2_2
timestamp 1743078376
transform 1 0 316 0 -1 105
box -2 -3 34 103
use BUFX2  BUFX2_5
timestamp 1743078376
transform -1 0 372 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_25
timestamp 1743078376
transform 1 0 316 0 1 105
box -2 -3 34 103
use INVX1  INVX1_16
timestamp 1743078376
transform -1 0 364 0 1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_7
timestamp 1743078376
transform 1 0 364 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_36
timestamp 1743078376
transform -1 0 404 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_13
timestamp 1743078376
transform -1 0 420 0 -1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_33
timestamp 1743078376
transform -1 0 452 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_31
timestamp 1743078376
transform -1 0 420 0 1 105
box -2 -3 34 103
use AND2X2  AND2X2_8
timestamp 1743078376
transform -1 0 452 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_28
timestamp 1743078376
transform -1 0 476 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_37
timestamp 1743078376
transform -1 0 508 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_23
timestamp 1743078376
transform -1 0 476 0 1 105
box -2 -3 26 103
use OAI22X1  OAI22X1_1
timestamp 1743078376
transform 1 0 476 0 1 105
box -2 -3 42 103
use NAND2X1  NAND2X1_14
timestamp 1743078376
transform 1 0 508 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_6
timestamp 1743078376
transform -1 0 548 0 -1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_13
timestamp 1743078376
transform -1 0 572 0 -1 105
box -2 -3 26 103
use AOI22X1  AOI22X1_7
timestamp 1743078376
transform -1 0 556 0 1 105
box -2 -3 42 103
use INVX4  INVX4_1
timestamp 1743078376
transform 1 0 572 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_1_0
timestamp 1743078376
transform 1 0 596 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1743078376
transform 1 0 604 0 -1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_4
timestamp 1743078376
transform 1 0 612 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_35
timestamp 1743078376
transform -1 0 588 0 1 105
box -2 -3 34 103
use AND2X2  AND2X2_7
timestamp 1743078376
transform 1 0 588 0 1 105
box -2 -3 34 103
use INVX1  INVX1_3
timestamp 1743078376
transform 1 0 636 0 -1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_40
timestamp 1743078376
transform 1 0 652 0 -1 105
box -2 -3 34 103
use FILL  FILL_1_1_0
timestamp 1743078376
transform 1 0 620 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_1
timestamp 1743078376
transform 1 0 628 0 1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_41
timestamp 1743078376
transform 1 0 636 0 1 105
box -2 -3 34 103
use AOI22X1  AOI22X1_8
timestamp 1743078376
transform 1 0 668 0 1 105
box -2 -3 42 103
use XNOR2X1  XNOR2X1_6
timestamp 1743078376
transform 1 0 684 0 -1 105
box -2 -3 58 103
use OR2X2  OR2X2_2
timestamp 1743078376
transform 1 0 708 0 1 105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_5
timestamp 1743078376
transform 1 0 740 0 -1 105
box -2 -3 58 103
use INVX1  INVX1_15
timestamp 1743078376
transform 1 0 796 0 -1 105
box -2 -3 18 103
use AOI21X1  AOI21X1_15
timestamp 1743078376
transform 1 0 740 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_3
timestamp 1743078376
transform 1 0 772 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_42
timestamp 1743078376
transform 1 0 812 0 -1 105
box -2 -3 34 103
use BUFX2  BUFX2_6
timestamp 1743078376
transform 1 0 844 0 -1 105
box -2 -3 26 103
use AND2X2  AND2X2_1
timestamp 1743078376
transform -1 0 836 0 1 105
box -2 -3 34 103
use INVX1  INVX1_4
timestamp 1743078376
transform -1 0 852 0 1 105
box -2 -3 18 103
use INVX2  INVX2_4
timestamp 1743078376
transform -1 0 868 0 1 105
box -2 -3 18 103
use FILL  FILL_1_1
timestamp 1743078376
transform -1 0 876 0 -1 105
box -2 -3 10 103
use FILL  FILL_2_1
timestamp 1743078376
transform 1 0 868 0 1 105
box -2 -3 10 103
use XOR2X1  XOR2X1_3
timestamp 1743078376
transform 1 0 4 0 -1 305
box -2 -3 58 103
use NAND2X1  NAND2X1_10
timestamp 1743078376
transform -1 0 84 0 -1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_3
timestamp 1743078376
transform 1 0 84 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_4
timestamp 1743078376
transform 1 0 116 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_21
timestamp 1743078376
transform 1 0 148 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_28
timestamp 1743078376
transform 1 0 172 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_24
timestamp 1743078376
transform 1 0 204 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_0_0
timestamp 1743078376
transform -1 0 244 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1743078376
transform -1 0 252 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_23
timestamp 1743078376
transform -1 0 284 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_8
timestamp 1743078376
transform 1 0 284 0 -1 305
box -2 -3 26 103
use INVX2  INVX2_7
timestamp 1743078376
transform -1 0 324 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_39
timestamp 1743078376
transform 1 0 324 0 -1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_6
timestamp 1743078376
transform -1 0 396 0 -1 305
box -2 -3 42 103
use NOR2X1  NOR2X1_25
timestamp 1743078376
transform 1 0 396 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_14
timestamp 1743078376
transform 1 0 420 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_34
timestamp 1743078376
transform 1 0 452 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_13
timestamp 1743078376
transform 1 0 484 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_14
timestamp 1743078376
transform 1 0 516 0 -1 305
box -2 -3 18 103
use OAI22X1  OAI22X1_2
timestamp 1743078376
transform -1 0 572 0 -1 305
box -2 -3 42 103
use NAND2X1  NAND2X1_15
timestamp 1743078376
transform 1 0 572 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_1_0
timestamp 1743078376
transform -1 0 604 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1743078376
transform -1 0 612 0 -1 305
box -2 -3 10 103
use NOR2X1  NOR2X1_11
timestamp 1743078376
transform -1 0 636 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_7
timestamp 1743078376
transform 1 0 636 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_16
timestamp 1743078376
transform -1 0 692 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_12
timestamp 1743078376
transform -1 0 716 0 -1 305
box -2 -3 26 103
use INVX4  INVX4_4
timestamp 1743078376
transform -1 0 740 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_7
timestamp 1743078376
transform 1 0 740 0 -1 305
box -2 -3 18 103
use AOI21X1  AOI21X1_5
timestamp 1743078376
transform 1 0 756 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_18
timestamp 1743078376
transform 1 0 788 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_45
timestamp 1743078376
transform 1 0 804 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_6
timestamp 1743078376
transform 1 0 836 0 -1 305
box -2 -3 26 103
use FILL  FILL_3_1
timestamp 1743078376
transform -1 0 868 0 -1 305
box -2 -3 10 103
use FILL  FILL_3_2
timestamp 1743078376
transform -1 0 876 0 -1 305
box -2 -3 10 103
use XNOR2X1  XNOR2X1_3
timestamp 1743078376
transform 1 0 4 0 1 305
box -2 -3 58 103
use OAI21X1  OAI21X1_21
timestamp 1743078376
transform -1 0 92 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_26
timestamp 1743078376
transform 1 0 92 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_43
timestamp 1743078376
transform 1 0 116 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_26
timestamp 1743078376
transform 1 0 148 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_27
timestamp 1743078376
transform 1 0 172 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_12
timestamp 1743078376
transform 1 0 204 0 1 305
box -2 -3 34 103
use FILL  FILL_3_0_0
timestamp 1743078376
transform -1 0 244 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1743078376
transform -1 0 252 0 1 305
box -2 -3 10 103
use INVX1  INVX1_12
timestamp 1743078376
transform -1 0 268 0 1 305
box -2 -3 18 103
use INVX1  INVX1_9
timestamp 1743078376
transform 1 0 268 0 1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_10
timestamp 1743078376
transform -1 0 308 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_27
timestamp 1743078376
transform -1 0 332 0 1 305
box -2 -3 26 103
use AOI22X1  AOI22X1_5
timestamp 1743078376
transform -1 0 372 0 1 305
box -2 -3 42 103
use AOI21X1  AOI21X1_7
timestamp 1743078376
transform 1 0 372 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_20
timestamp 1743078376
transform 1 0 404 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_8
timestamp 1743078376
transform 1 0 428 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_16
timestamp 1743078376
transform 1 0 460 0 1 305
box -2 -3 34 103
use INVX1  INVX1_17
timestamp 1743078376
transform -1 0 508 0 1 305
box -2 -3 18 103
use AOI21X1  AOI21X1_8
timestamp 1743078376
transform 1 0 508 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_48
timestamp 1743078376
transform -1 0 572 0 1 305
box -2 -3 34 103
use INVX2  INVX2_13
timestamp 1743078376
transform 1 0 572 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_44
timestamp 1743078376
transform 1 0 588 0 1 305
box -2 -3 34 103
use FILL  FILL_3_1_0
timestamp 1743078376
transform 1 0 620 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1743078376
transform 1 0 628 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_49
timestamp 1743078376
transform 1 0 636 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_27
timestamp 1743078376
transform -1 0 692 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_9
timestamp 1743078376
transform 1 0 692 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_29
timestamp 1743078376
transform 1 0 724 0 1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_5
timestamp 1743078376
transform -1 0 780 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_6
timestamp 1743078376
transform 1 0 780 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_46
timestamp 1743078376
transform 1 0 812 0 1 305
box -2 -3 34 103
use BUFX2  BUFX2_7
timestamp 1743078376
transform 1 0 844 0 1 305
box -2 -3 26 103
use FILL  FILL_4_1
timestamp 1743078376
transform 1 0 868 0 1 305
box -2 -3 10 103
use BUFX2  BUFX2_2
timestamp 1743078376
transform -1 0 28 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_3
timestamp 1743078376
transform -1 0 60 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_20
timestamp 1743078376
transform -1 0 92 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_15
timestamp 1743078376
transform -1 0 124 0 -1 505
box -2 -3 34 103
use AND2X2  AND2X2_5
timestamp 1743078376
transform -1 0 156 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_19
timestamp 1743078376
transform 1 0 156 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_10
timestamp 1743078376
transform -1 0 220 0 -1 505
box -2 -3 34 103
use INVX2  INVX2_11
timestamp 1743078376
transform -1 0 236 0 -1 505
box -2 -3 18 103
use FILL  FILL_4_0_0
timestamp 1743078376
transform 1 0 236 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1743078376
transform 1 0 244 0 -1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_17
timestamp 1743078376
transform 1 0 252 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_19
timestamp 1743078376
transform 1 0 284 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_18
timestamp 1743078376
transform 1 0 308 0 -1 505
box -2 -3 34 103
use AOI22X1  AOI22X1_4
timestamp 1743078376
transform -1 0 380 0 -1 505
box -2 -3 42 103
use INVX4  INVX4_3
timestamp 1743078376
transform -1 0 404 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_15
timestamp 1743078376
transform 1 0 404 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_10
timestamp 1743078376
transform -1 0 460 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_2
timestamp 1743078376
transform 1 0 460 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_18
timestamp 1743078376
transform -1 0 508 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_16
timestamp 1743078376
transform 1 0 508 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_47
timestamp 1743078376
transform -1 0 564 0 -1 505
box -2 -3 34 103
use INVX2  INVX2_12
timestamp 1743078376
transform -1 0 580 0 -1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_18
timestamp 1743078376
transform -1 0 604 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_1_0
timestamp 1743078376
transform 1 0 604 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1743078376
transform 1 0 612 0 -1 505
box -2 -3 10 103
use NAND2X1  NAND2X1_1
timestamp 1743078376
transform 1 0 620 0 -1 505
box -2 -3 26 103
use AOI22X1  AOI22X1_9
timestamp 1743078376
transform -1 0 684 0 -1 505
box -2 -3 42 103
use INVX4  INVX4_2
timestamp 1743078376
transform -1 0 708 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_21
timestamp 1743078376
transform -1 0 732 0 -1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_7
timestamp 1743078376
transform -1 0 764 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_8
timestamp 1743078376
transform -1 0 796 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_2
timestamp 1743078376
transform 1 0 796 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_17
timestamp 1743078376
transform -1 0 852 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_30
timestamp 1743078376
transform -1 0 876 0 -1 505
box -2 -3 26 103
use INVX2  INVX2_5
timestamp 1743078376
transform 1 0 4 0 1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_6
timestamp 1743078376
transform 1 0 20 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_8
timestamp 1743078376
transform -1 0 68 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_9
timestamp 1743078376
transform -1 0 100 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_9
timestamp 1743078376
transform -1 0 124 0 1 505
box -2 -3 26 103
use INVX1  INVX1_8
timestamp 1743078376
transform 1 0 124 0 1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_25
timestamp 1743078376
transform -1 0 164 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_38
timestamp 1743078376
transform -1 0 196 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_6
timestamp 1743078376
transform -1 0 228 0 1 505
box -2 -3 34 103
use FILL  FILL_5_0_0
timestamp 1743078376
transform 1 0 228 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1743078376
transform 1 0 236 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_16
timestamp 1743078376
transform 1 0 244 0 1 505
box -2 -3 34 103
use XOR2X1  XOR2X1_1
timestamp 1743078376
transform 1 0 276 0 1 505
box -2 -3 58 103
use AOI22X1  AOI22X1_3
timestamp 1743078376
transform -1 0 372 0 1 505
box -2 -3 42 103
use NAND2X1  NAND2X1_24
timestamp 1743078376
transform 1 0 372 0 1 505
box -2 -3 26 103
use INVX1  INVX1_11
timestamp 1743078376
transform -1 0 412 0 1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_23
timestamp 1743078376
transform 1 0 412 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_3
timestamp 1743078376
transform 1 0 436 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_13
timestamp 1743078376
transform 1 0 460 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_14
timestamp 1743078376
transform -1 0 508 0 1 505
box -2 -3 26 103
use INVX2  INVX2_2
timestamp 1743078376
transform 1 0 508 0 1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_4
timestamp 1743078376
transform 1 0 524 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_3
timestamp 1743078376
transform -1 0 572 0 1 505
box -2 -3 26 103
use INVX2  INVX2_3
timestamp 1743078376
transform 1 0 572 0 1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_5
timestamp 1743078376
transform 1 0 588 0 1 505
box -2 -3 26 103
use FILL  FILL_5_1_0
timestamp 1743078376
transform 1 0 612 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1743078376
transform 1 0 620 0 1 505
box -2 -3 10 103
use NAND3X1  NAND3X1_2
timestamp 1743078376
transform 1 0 628 0 1 505
box -2 -3 34 103
use AOI22X1  AOI22X1_1
timestamp 1743078376
transform 1 0 660 0 1 505
box -2 -3 42 103
use INVX2  INVX2_8
timestamp 1743078376
transform -1 0 716 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_5
timestamp 1743078376
transform -1 0 748 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_1
timestamp 1743078376
transform 1 0 748 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_2
timestamp 1743078376
transform -1 0 812 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_1
timestamp 1743078376
transform 1 0 812 0 1 505
box -2 -3 34 103
use BUFX2  BUFX2_8
timestamp 1743078376
transform 1 0 844 0 1 505
box -2 -3 26 103
use FILL  FILL_6_1
timestamp 1743078376
transform 1 0 868 0 1 505
box -2 -3 10 103
use NAND2X1  NAND2X1_9
timestamp 1743078376
transform 1 0 4 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_5
timestamp 1743078376
transform -1 0 44 0 -1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_19
timestamp 1743078376
transform 1 0 44 0 -1 705
box -2 -3 26 103
use INVX2  INVX2_9
timestamp 1743078376
transform 1 0 68 0 -1 705
box -2 -3 18 103
use INVX1  INVX1_10
timestamp 1743078376
transform 1 0 84 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_11
timestamp 1743078376
transform 1 0 100 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_24
timestamp 1743078376
transform -1 0 156 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_13
timestamp 1743078376
transform 1 0 156 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_12
timestamp 1743078376
transform -1 0 220 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_17
timestamp 1743078376
transform 1 0 220 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_0_0
timestamp 1743078376
transform 1 0 244 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1743078376
transform 1 0 252 0 -1 705
box -2 -3 10 103
use AND2X2  AND2X2_4
timestamp 1743078376
transform 1 0 260 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_22
timestamp 1743078376
transform 1 0 292 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_1
timestamp 1743078376
transform -1 0 340 0 -1 705
box -2 -3 26 103
use INVX2  INVX2_1
timestamp 1743078376
transform 1 0 340 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_2
timestamp 1743078376
transform 1 0 356 0 -1 705
box -2 -3 34 103
use OR2X2  OR2X2_1
timestamp 1743078376
transform 1 0 388 0 -1 705
box -2 -3 34 103
use INVX2  INVX2_10
timestamp 1743078376
transform 1 0 420 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_14
timestamp 1743078376
transform -1 0 468 0 -1 705
box -2 -3 34 103
use BUFX2  BUFX2_1
timestamp 1743078376
transform 1 0 468 0 -1 705
box -2 -3 26 103
use AOI22X1  AOI22X1_2
timestamp 1743078376
transform -1 0 532 0 -1 705
box -2 -3 42 103
use NOR2X1  NOR2X1_12
timestamp 1743078376
transform -1 0 556 0 -1 705
box -2 -3 26 103
use AND2X2  AND2X2_3
timestamp 1743078376
transform -1 0 588 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_1
timestamp 1743078376
transform 1 0 588 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_1_0
timestamp 1743078376
transform 1 0 620 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1743078376
transform 1 0 628 0 -1 705
box -2 -3 10 103
use INVX1  INVX1_1
timestamp 1743078376
transform 1 0 636 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_6
timestamp 1743078376
transform 1 0 652 0 -1 705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_1
timestamp 1743078376
transform 1 0 684 0 -1 705
box -2 -3 58 103
use NAND2X1  NAND2X1_17
timestamp 1743078376
transform -1 0 764 0 -1 705
box -2 -3 26 103
use BUFX2  BUFX2_9
timestamp 1743078376
transform 1 0 764 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_5
timestamp 1743078376
transform 1 0 788 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_7
timestamp 1743078376
transform 1 0 812 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_2
timestamp 1743078376
transform -1 0 852 0 -1 705
box -2 -3 18 103
use FILL  FILL_7_1
timestamp 1743078376
transform -1 0 860 0 -1 705
box -2 -3 10 103
use FILL  FILL_7_2
timestamp 1743078376
transform -1 0 868 0 -1 705
box -2 -3 10 103
use FILL  FILL_7_3
timestamp 1743078376
transform -1 0 876 0 -1 705
box -2 -3 10 103
<< labels >>
flabel metal6 s 232 -30 248 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 608 -30 624 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 150 728 154 732 3 FreeSans 24 90 0 0 A[0]
port 2 nsew
flabel metal3 s -26 548 -22 552 7 FreeSans 24 0 0 0 A[1]
port 3 nsew
flabel metal3 s -26 268 -22 272 7 FreeSans 24 0 0 0 A[2]
port 4 nsew
flabel metal2 s 302 -22 306 -18 7 FreeSans 24 270 0 0 A[3]
port 5 nsew
flabel metal2 s 574 -22 578 -18 7 FreeSans 24 270 0 0 A[4]
port 6 nsew
flabel metal3 s 902 148 906 152 3 FreeSans 24 0 0 0 A[5]
port 7 nsew
flabel metal2 s 510 728 514 732 3 FreeSans 24 90 0 0 A[6]
port 8 nsew
flabel metal2 s 630 728 634 732 3 FreeSans 24 90 0 0 A[7]
port 9 nsew
flabel metal3 s -26 648 -22 652 7 FreeSans 24 90 0 0 B[0]
port 10 nsew
flabel metal3 s -26 528 -22 532 7 FreeSans 24 0 0 0 B[1]
port 11 nsew
flabel metal3 s -26 288 -22 292 7 FreeSans 24 0 0 0 B[2]
port 12 nsew
flabel metal2 s 326 -22 330 -18 7 FreeSans 24 270 0 0 B[3]
port 13 nsew
flabel metal2 s 550 -22 554 -18 7 FreeSans 24 270 0 0 B[4]
port 14 nsew
flabel metal3 s 902 558 906 562 3 FreeSans 24 0 0 0 B[5]
port 15 nsew
flabel metal2 s 534 728 538 732 3 FreeSans 24 90 0 0 B[6]
port 16 nsew
flabel metal2 s 710 728 714 732 3 FreeSans 24 90 0 0 B[7]
port 17 nsew
flabel metal2 s 302 728 306 732 3 FreeSans 24 90 0 0 ALU_Sel[0]
port 18 nsew
flabel metal2 s 326 728 330 732 3 FreeSans 24 90 0 0 ALU_Sel[1]
port 19 nsew
flabel metal2 s 222 728 226 732 3 FreeSans 24 90 0 0 ALU_Sel[2]
port 20 nsew
flabel metal2 s 478 728 482 732 3 FreeSans 24 90 0 0 ALU_Out[0]
port 21 nsew
flabel metal3 s -26 448 -22 452 7 FreeSans 24 0 0 0 ALU_Out[1]
port 22 nsew
flabel metal3 s -26 148 -22 152 7 FreeSans 24 0 0 0 ALU_Out[2]
port 23 nsew
flabel metal3 s -26 48 -22 52 7 FreeSans 24 270 0 0 ALU_Out[3]
port 24 nsew
flabel metal2 s 358 -22 362 -18 7 FreeSans 24 270 0 0 ALU_Out[4]
port 25 nsew
flabel metal2 s 854 -22 858 -18 3 FreeSans 24 270 0 0 ALU_Out[5]
port 26 nsew
flabel metal3 s 902 348 906 352 3 FreeSans 24 0 0 0 ALU_Out[6]
port 27 nsew
flabel metal3 s 902 578 906 582 3 FreeSans 24 0 0 0 ALU_Out[7]
port 28 nsew
flabel metal2 s 774 728 778 732 3 FreeSans 24 90 0 0 CarryOut
port 29 nsew
<< end >>
