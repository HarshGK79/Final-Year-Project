VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ALU_8bit
  CLASS BLOCK ;
  FOREIGN ALU_8bit ;
  ORIGIN 2.600 3.000 ;
  SIZE 93.200 BY 76.200 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.600 60.800 1.000 63.100 ;
        RECT 2.200 60.800 2.600 63.100 ;
        RECT 3.800 60.800 4.200 63.100 ;
        RECT 4.600 60.800 5.000 63.100 ;
        RECT 6.200 60.800 6.600 63.100 ;
        RECT 7.000 60.800 7.400 65.100 ;
        RECT 8.600 60.800 9.000 63.100 ;
        RECT 10.200 60.800 10.600 65.100 ;
        RECT 12.300 60.800 12.700 63.100 ;
        RECT 15.000 60.800 15.400 65.100 ;
        RECT 15.800 60.800 16.200 65.100 ;
        RECT 17.900 60.800 18.300 63.100 ;
        RECT 19.300 60.800 19.700 63.100 ;
        RECT 21.400 60.800 21.800 65.100 ;
        RECT 22.200 60.800 22.600 65.100 ;
        RECT 26.200 60.800 26.600 63.100 ;
        RECT 27.800 60.800 28.200 64.900 ;
        RECT 29.400 60.800 29.800 63.100 ;
        RECT 31.000 60.800 31.400 63.100 ;
        RECT 33.400 60.800 33.800 65.100 ;
        RECT 34.200 60.800 34.600 65.100 ;
        RECT 35.800 60.800 36.200 65.100 ;
        RECT 37.900 60.800 38.300 63.100 ;
        RECT 40.300 60.800 40.700 65.100 ;
        RECT 42.200 60.800 42.600 65.100 ;
        RECT 44.100 60.800 44.500 63.100 ;
        RECT 46.200 60.800 46.600 65.100 ;
        RECT 47.800 60.800 48.200 64.500 ;
        RECT 51.800 60.800 52.200 64.500 ;
        RECT 55.000 60.800 55.400 65.100 ;
        RECT 56.600 60.800 57.000 64.900 ;
        RECT 58.200 60.800 58.600 63.100 ;
        RECT 59.000 60.800 59.400 65.100 ;
        RECT 61.100 60.800 61.500 63.100 ;
        RECT 63.800 60.800 64.200 63.100 ;
        RECT 65.400 60.800 65.800 65.100 ;
        RECT 67.500 60.800 67.900 63.100 ;
        RECT 69.400 61.100 69.900 64.400 ;
        RECT 69.500 60.800 69.900 61.100 ;
        RECT 72.500 60.800 73.000 64.400 ;
        RECT 74.200 60.800 74.600 63.100 ;
        RECT 75.800 60.800 76.200 63.100 ;
        RECT 77.400 60.800 77.800 64.500 ;
        RECT 79.000 60.800 79.400 65.100 ;
        RECT 81.400 60.800 81.800 63.100 ;
        RECT 83.000 60.800 83.400 63.100 ;
        RECT 84.600 60.800 85.000 63.100 ;
        RECT 0.200 60.200 87.800 60.800 ;
        RECT 0.600 55.900 1.000 60.200 ;
        RECT 2.200 55.900 2.600 60.200 ;
        RECT 4.600 57.900 5.000 60.200 ;
        RECT 6.200 57.900 6.600 60.200 ;
        RECT 8.600 56.500 9.000 60.200 ;
        RECT 11.800 55.900 12.200 60.200 ;
        RECT 12.600 57.900 13.000 60.200 ;
        RECT 14.200 57.900 14.600 60.200 ;
        RECT 15.800 57.900 16.200 60.200 ;
        RECT 16.900 57.900 17.300 60.200 ;
        RECT 19.000 55.900 19.400 60.200 ;
        RECT 21.400 56.500 21.800 60.200 ;
        RECT 24.600 55.900 25.000 60.200 ;
        RECT 26.700 57.900 27.100 60.200 ;
        RECT 28.700 59.900 29.100 60.200 ;
        RECT 28.600 56.600 29.100 59.900 ;
        RECT 31.700 56.600 32.200 60.200 ;
        RECT 35.800 56.500 36.200 60.200 ;
        RECT 37.400 57.900 37.800 60.200 ;
        RECT 39.000 57.900 39.400 60.200 ;
        RECT 40.600 57.900 41.000 60.200 ;
        RECT 41.400 57.900 41.800 60.200 ;
        RECT 43.000 57.900 43.400 60.200 ;
        RECT 43.800 57.900 44.200 60.200 ;
        RECT 45.400 57.900 45.800 60.200 ;
        RECT 46.200 55.900 46.600 60.200 ;
        RECT 50.200 55.900 50.600 60.200 ;
        RECT 51.000 55.900 51.400 60.200 ;
        RECT 52.600 57.900 53.000 60.200 ;
        RECT 54.200 57.900 54.600 60.200 ;
        RECT 56.600 55.900 57.000 60.200 ;
        RECT 57.400 55.900 57.800 60.200 ;
        RECT 59.000 57.900 59.400 60.200 ;
        RECT 60.600 57.900 61.000 60.200 ;
        RECT 63.000 57.900 63.400 60.200 ;
        RECT 64.600 58.100 65.000 60.200 ;
        RECT 67.000 56.500 67.400 60.200 ;
        RECT 71.000 55.900 71.400 60.200 ;
        RECT 72.100 57.900 72.500 60.200 ;
        RECT 74.200 55.900 74.600 60.200 ;
        RECT 75.800 56.500 76.200 60.200 ;
        RECT 79.800 56.500 80.200 60.200 ;
        RECT 81.400 57.900 81.800 60.200 ;
        RECT 83.000 58.100 83.400 60.200 ;
        RECT 85.400 56.500 85.800 60.200 ;
        RECT 1.400 40.800 1.800 44.500 ;
        RECT 4.600 40.800 5.000 44.500 ;
        RECT 6.500 40.800 6.900 43.100 ;
        RECT 8.600 40.800 9.000 45.100 ;
        RECT 9.700 40.800 10.100 43.100 ;
        RECT 11.800 40.800 12.200 45.100 ;
        RECT 13.400 40.800 13.800 44.900 ;
        RECT 15.000 40.800 15.400 43.100 ;
        RECT 15.800 40.800 16.200 45.100 ;
        RECT 17.900 40.800 18.300 43.100 ;
        RECT 20.600 40.800 21.000 44.500 ;
        RECT 23.000 40.800 23.400 45.100 ;
        RECT 25.400 40.800 25.800 45.100 ;
        RECT 27.500 40.800 27.900 43.100 ;
        RECT 28.600 40.800 29.000 45.100 ;
        RECT 31.000 40.800 31.400 45.100 ;
        RECT 33.100 40.800 33.500 43.100 ;
        RECT 36.600 40.800 37.000 44.500 ;
        RECT 38.200 40.800 38.600 45.100 ;
        RECT 39.800 40.800 40.200 45.100 ;
        RECT 40.600 40.800 41.000 45.100 ;
        RECT 43.300 40.800 43.700 43.100 ;
        RECT 45.400 40.800 45.800 45.100 ;
        RECT 46.200 40.800 46.600 45.100 ;
        RECT 50.200 40.800 50.600 45.100 ;
        RECT 51.000 40.800 51.400 45.100 ;
        RECT 53.700 40.800 54.100 43.100 ;
        RECT 55.800 40.800 56.200 45.100 ;
        RECT 57.400 40.800 57.800 45.100 ;
        RECT 58.200 40.800 58.600 43.100 ;
        RECT 59.800 40.800 60.200 43.100 ;
        RECT 62.200 40.800 62.600 43.100 ;
        RECT 63.800 40.800 64.200 43.100 ;
        RECT 67.000 40.800 67.400 44.500 ;
        RECT 68.600 40.800 69.000 45.100 ;
        RECT 70.200 40.800 70.600 45.100 ;
        RECT 71.000 40.800 71.400 43.100 ;
        RECT 72.600 40.800 73.000 43.100 ;
        RECT 74.200 40.800 74.600 42.900 ;
        RECT 75.800 40.800 76.200 43.100 ;
        RECT 77.400 40.800 77.800 42.900 ;
        RECT 79.000 40.800 79.400 43.100 ;
        RECT 79.800 40.800 80.200 43.100 ;
        RECT 81.400 40.800 81.800 43.100 ;
        RECT 83.800 40.800 84.200 44.500 ;
        RECT 85.400 40.800 85.800 43.100 ;
        RECT 87.000 40.800 87.400 43.100 ;
        RECT 0.200 40.200 87.800 40.800 ;
        RECT 1.500 39.900 1.900 40.200 ;
        RECT 1.400 36.600 1.900 39.900 ;
        RECT 4.500 36.600 5.000 40.200 ;
        RECT 6.500 37.900 6.900 40.200 ;
        RECT 8.600 35.900 9.000 40.200 ;
        RECT 9.400 37.900 9.800 40.200 ;
        RECT 11.000 37.900 11.400 40.200 ;
        RECT 11.800 35.900 12.200 40.200 ;
        RECT 13.900 37.900 14.300 40.200 ;
        RECT 15.000 35.900 15.400 40.200 ;
        RECT 17.400 35.900 17.800 40.200 ;
        RECT 19.500 37.900 19.900 40.200 ;
        RECT 21.400 36.500 21.800 40.200 ;
        RECT 26.200 37.900 26.600 40.200 ;
        RECT 27.000 37.900 27.400 40.200 ;
        RECT 30.200 35.900 30.600 40.200 ;
        RECT 31.000 37.900 31.400 40.200 ;
        RECT 32.600 37.900 33.000 40.200 ;
        RECT 35.800 36.500 36.200 40.200 ;
        RECT 38.200 36.500 38.600 40.200 ;
        RECT 40.600 37.900 41.000 40.200 ;
        RECT 42.200 37.900 42.600 40.200 ;
        RECT 43.000 35.900 43.400 40.200 ;
        RECT 45.100 37.900 45.500 40.200 ;
        RECT 47.000 36.500 47.400 40.200 ;
        RECT 50.200 37.900 50.600 40.200 ;
        RECT 51.800 36.500 52.200 40.200 ;
        RECT 54.500 37.900 54.900 40.200 ;
        RECT 56.600 35.900 57.000 40.200 ;
        RECT 57.400 35.900 57.800 40.200 ;
        RECT 59.000 35.900 59.400 40.200 ;
        RECT 61.100 37.900 61.500 40.200 ;
        RECT 63.800 35.900 64.200 40.200 ;
        RECT 65.900 37.900 66.300 40.200 ;
        RECT 68.600 35.900 69.000 40.200 ;
        RECT 69.400 35.900 69.800 40.200 ;
        RECT 71.500 37.900 71.900 40.200 ;
        RECT 72.600 37.900 73.000 40.200 ;
        RECT 74.200 37.900 74.600 40.200 ;
        RECT 75.800 38.100 76.200 40.200 ;
        RECT 77.400 37.900 77.800 40.200 ;
        RECT 78.200 37.900 78.600 40.200 ;
        RECT 79.800 38.100 80.200 40.200 ;
        RECT 81.400 35.900 81.800 40.200 ;
        RECT 83.500 37.900 83.900 40.200 ;
        RECT 85.400 36.500 85.800 40.200 ;
        RECT 1.400 21.100 1.900 24.400 ;
        RECT 1.500 20.800 1.900 21.100 ;
        RECT 4.500 20.800 5.000 24.400 ;
        RECT 6.200 20.800 6.600 23.100 ;
        RECT 7.800 20.800 8.200 23.100 ;
        RECT 8.600 20.800 9.000 23.100 ;
        RECT 10.200 20.800 10.600 22.900 ;
        RECT 11.800 20.800 12.200 25.100 ;
        RECT 13.900 20.800 14.300 23.100 ;
        RECT 15.000 20.800 15.400 25.100 ;
        RECT 17.400 20.800 17.800 25.100 ;
        RECT 19.500 20.800 19.900 23.100 ;
        RECT 20.600 20.800 21.000 25.100 ;
        RECT 22.700 20.800 23.100 23.100 ;
        RECT 25.700 20.800 26.100 23.100 ;
        RECT 27.800 20.800 28.200 25.100 ;
        RECT 28.600 20.800 29.000 25.100 ;
        RECT 31.800 20.800 32.200 25.100 ;
        RECT 32.600 20.800 33.000 25.100 ;
        RECT 34.700 20.800 35.100 23.100 ;
        RECT 38.200 20.800 38.600 24.500 ;
        RECT 39.800 20.800 40.200 25.100 ;
        RECT 43.000 20.800 43.400 24.500 ;
        RECT 45.400 20.800 45.800 25.100 ;
        RECT 47.500 20.800 47.900 23.100 ;
        RECT 49.400 20.800 49.800 24.500 ;
        RECT 51.800 20.800 52.200 23.100 ;
        RECT 53.400 20.800 53.800 25.100 ;
        RECT 56.600 20.800 57.000 25.100 ;
        RECT 57.400 20.800 57.800 23.100 ;
        RECT 59.000 20.800 59.400 23.100 ;
        RECT 63.000 20.800 63.400 25.100 ;
        RECT 63.800 20.800 64.200 25.100 ;
        RECT 65.900 20.800 66.300 23.100 ;
        RECT 67.000 20.800 67.400 23.100 ;
        RECT 68.600 20.800 69.000 23.100 ;
        RECT 69.400 20.800 69.800 23.100 ;
        RECT 71.000 20.800 71.400 23.100 ;
        RECT 71.800 20.800 72.200 25.100 ;
        RECT 73.400 20.800 73.800 25.100 ;
        RECT 74.200 20.800 74.600 23.100 ;
        RECT 76.600 20.800 77.000 24.500 ;
        RECT 79.000 20.800 79.400 23.100 ;
        RECT 80.600 20.800 81.000 25.100 ;
        RECT 82.700 20.800 83.100 23.100 ;
        RECT 83.800 20.800 84.200 23.100 ;
        RECT 85.400 20.800 85.800 23.100 ;
        RECT 0.200 20.200 87.800 20.800 ;
        RECT 1.400 16.500 1.800 20.200 ;
        RECT 3.800 18.100 4.200 20.200 ;
        RECT 5.400 17.900 5.800 20.200 ;
        RECT 6.200 15.900 6.600 20.200 ;
        RECT 8.300 17.900 8.700 20.200 ;
        RECT 11.000 16.500 11.400 20.200 ;
        RECT 12.600 15.900 13.000 20.200 ;
        RECT 14.700 17.900 15.100 20.200 ;
        RECT 17.400 15.900 17.800 20.200 ;
        RECT 18.200 15.900 18.600 20.200 ;
        RECT 20.300 17.900 20.700 20.200 ;
        RECT 21.400 15.900 21.800 20.200 ;
        RECT 25.700 17.900 26.100 20.200 ;
        RECT 27.800 15.900 28.200 20.200 ;
        RECT 29.400 16.500 29.800 20.200 ;
        RECT 31.800 15.900 32.200 20.200 ;
        RECT 33.900 17.900 34.300 20.200 ;
        RECT 35.800 17.900 36.200 20.200 ;
        RECT 36.600 15.900 37.000 20.200 ;
        RECT 39.300 17.900 39.700 20.200 ;
        RECT 41.400 15.900 41.800 20.200 ;
        RECT 43.000 16.100 43.400 20.200 ;
        RECT 44.600 17.900 45.000 20.200 ;
        RECT 47.000 15.900 47.400 20.200 ;
        RECT 47.800 15.900 48.200 20.200 ;
        RECT 51.000 15.900 51.400 20.200 ;
        RECT 54.200 16.500 54.600 20.200 ;
        RECT 56.100 17.900 56.500 20.200 ;
        RECT 58.200 15.900 58.600 20.200 ;
        RECT 59.000 17.900 59.400 20.200 ;
        RECT 60.600 16.100 61.000 20.200 ;
        RECT 63.800 15.900 64.200 20.200 ;
        RECT 65.900 17.900 66.300 20.200 ;
        RECT 67.800 16.500 68.200 20.200 ;
        RECT 72.300 15.900 72.700 20.200 ;
        RECT 75.000 16.500 75.400 20.200 ;
        RECT 77.400 15.900 77.800 20.200 ;
        RECT 79.500 17.900 79.900 20.200 ;
        RECT 81.400 16.100 81.800 20.200 ;
        RECT 83.000 17.900 83.400 20.200 ;
        RECT 84.600 17.900 85.000 20.200 ;
        RECT 86.200 15.900 86.600 20.200 ;
        RECT 1.400 0.800 1.800 4.500 ;
        RECT 3.800 1.100 4.300 4.400 ;
        RECT 3.900 0.800 4.300 1.100 ;
        RECT 6.900 0.800 7.400 4.400 ;
        RECT 8.600 0.800 9.000 5.100 ;
        RECT 10.700 0.800 11.100 3.100 ;
        RECT 12.600 0.800 13.000 4.900 ;
        RECT 14.200 0.800 14.600 3.100 ;
        RECT 15.800 1.100 16.300 4.400 ;
        RECT 15.900 0.800 16.300 1.100 ;
        RECT 18.900 0.800 19.400 4.400 ;
        RECT 21.400 0.800 21.900 4.400 ;
        RECT 24.500 1.100 25.000 4.400 ;
        RECT 24.500 0.800 24.900 1.100 ;
        RECT 27.800 0.800 28.200 3.100 ;
        RECT 29.400 0.800 29.800 3.100 ;
        RECT 30.200 0.800 30.600 5.100 ;
        RECT 31.800 0.800 32.200 3.100 ;
        RECT 33.400 0.800 33.800 4.900 ;
        RECT 35.800 0.800 36.200 4.500 ;
        RECT 37.700 0.800 38.100 3.100 ;
        RECT 39.800 0.800 40.200 5.100 ;
        RECT 41.400 0.800 41.800 3.100 ;
        RECT 42.500 0.800 42.900 3.100 ;
        RECT 44.600 0.800 45.000 5.100 ;
        RECT 45.400 0.800 45.800 3.100 ;
        RECT 47.000 0.800 47.400 3.100 ;
        RECT 48.100 0.800 48.500 3.100 ;
        RECT 50.200 0.800 50.600 5.100 ;
        RECT 51.000 0.800 51.400 3.100 ;
        RECT 52.600 0.800 53.000 3.100 ;
        RECT 54.200 0.800 54.600 3.100 ;
        RECT 55.000 0.800 55.400 3.100 ;
        RECT 56.600 0.800 57.000 3.100 ;
        RECT 57.400 0.800 57.800 5.100 ;
        RECT 59.000 0.800 59.400 5.100 ;
        RECT 61.400 0.800 61.800 5.100 ;
        RECT 63.800 0.800 64.200 3.100 ;
        RECT 65.400 0.800 65.800 5.100 ;
        RECT 67.500 0.800 67.900 3.100 ;
        RECT 69.400 1.100 69.900 4.400 ;
        RECT 69.500 0.800 69.900 1.100 ;
        RECT 72.500 0.800 73.000 4.400 ;
        RECT 75.000 1.100 75.500 4.400 ;
        RECT 75.100 0.800 75.500 1.100 ;
        RECT 78.100 0.800 78.600 4.400 ;
        RECT 79.800 0.800 80.200 3.100 ;
        RECT 81.400 0.800 81.800 5.100 ;
        RECT 83.500 0.800 83.900 3.100 ;
        RECT 85.400 0.800 85.800 4.500 ;
        RECT 0.200 0.200 87.800 0.800 ;
      LAYER via1 ;
        RECT 23.400 60.300 23.800 60.700 ;
        RECT 24.100 60.300 24.500 60.700 ;
        RECT 23.400 40.300 23.800 40.700 ;
        RECT 24.100 40.300 24.500 40.700 ;
        RECT 23.400 20.300 23.800 20.700 ;
        RECT 24.100 20.300 24.500 20.700 ;
        RECT 23.400 0.300 23.800 0.700 ;
        RECT 24.100 0.300 24.500 0.700 ;
      LAYER metal2 ;
        RECT 23.200 60.300 24.800 60.700 ;
        RECT 23.200 40.300 24.800 40.700 ;
        RECT 23.200 20.300 24.800 20.700 ;
        RECT 23.200 0.300 24.800 0.700 ;
      LAYER via2 ;
        RECT 23.400 60.300 23.800 60.700 ;
        RECT 24.100 60.300 24.500 60.700 ;
        RECT 23.400 40.300 23.800 40.700 ;
        RECT 24.100 40.300 24.500 40.700 ;
        RECT 23.400 20.300 23.800 20.700 ;
        RECT 24.100 20.300 24.500 20.700 ;
        RECT 23.400 0.300 23.800 0.700 ;
        RECT 24.100 0.300 24.500 0.700 ;
      LAYER metal3 ;
        RECT 23.200 60.300 24.800 60.700 ;
        RECT 23.200 40.300 24.800 40.700 ;
        RECT 23.200 20.300 24.800 20.700 ;
        RECT 23.200 0.300 24.800 0.700 ;
      LAYER via3 ;
        RECT 23.400 60.300 23.800 60.700 ;
        RECT 24.200 60.300 24.600 60.700 ;
        RECT 23.400 40.300 23.800 40.700 ;
        RECT 24.200 40.300 24.600 40.700 ;
        RECT 23.400 20.300 23.800 20.700 ;
        RECT 24.200 20.300 24.600 20.700 ;
        RECT 23.400 0.300 23.800 0.700 ;
        RECT 24.200 0.300 24.600 0.700 ;
      LAYER metal4 ;
        RECT 23.200 60.300 24.800 60.700 ;
        RECT 23.200 40.300 24.800 40.700 ;
        RECT 23.200 20.300 24.800 20.700 ;
        RECT 23.200 0.300 24.800 0.700 ;
      LAYER via4 ;
        RECT 23.400 60.300 23.800 60.700 ;
        RECT 24.100 60.300 24.500 60.700 ;
        RECT 23.400 40.300 23.800 40.700 ;
        RECT 24.100 40.300 24.500 40.700 ;
        RECT 23.400 20.300 23.800 20.700 ;
        RECT 24.100 20.300 24.500 20.700 ;
        RECT 23.400 0.300 23.800 0.700 ;
        RECT 24.100 0.300 24.500 0.700 ;
      LAYER metal5 ;
        RECT 23.200 60.200 24.800 60.700 ;
        RECT 23.200 40.200 24.800 40.700 ;
        RECT 23.200 20.200 24.800 20.700 ;
        RECT 23.200 0.200 24.800 0.700 ;
      LAYER via5 ;
        RECT 24.200 60.200 24.700 60.700 ;
        RECT 24.200 40.200 24.700 40.700 ;
        RECT 24.200 20.200 24.700 20.700 ;
        RECT 24.200 0.200 24.700 0.700 ;
      LAYER metal6 ;
        RECT 23.200 -3.000 24.800 73.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.200 70.200 87.800 70.800 ;
        RECT 0.600 67.900 1.000 70.200 ;
        RECT 3.800 68.900 4.200 70.200 ;
        RECT 4.600 67.900 5.000 70.200 ;
        RECT 7.000 67.900 7.400 70.200 ;
        RECT 8.600 68.900 9.000 70.200 ;
        RECT 11.000 68.300 11.400 70.200 ;
        RECT 13.400 68.900 13.800 70.200 ;
        RECT 15.000 68.900 15.400 70.200 ;
        RECT 16.600 68.300 17.000 70.200 ;
        RECT 20.600 68.300 21.000 70.200 ;
        RECT 22.200 68.900 22.600 70.200 ;
        RECT 23.800 68.900 24.200 70.200 ;
        RECT 27.500 68.000 27.900 70.200 ;
        RECT 29.400 67.900 29.800 70.200 ;
        RECT 31.800 68.900 32.200 70.200 ;
        RECT 33.400 68.900 33.800 70.200 ;
        RECT 34.200 67.900 34.600 70.200 ;
        RECT 36.600 68.300 37.000 70.200 ;
        RECT 39.000 68.900 39.400 70.200 ;
        RECT 40.600 68.100 41.000 70.200 ;
        RECT 42.200 67.900 42.600 70.200 ;
        RECT 45.400 68.300 45.800 70.200 ;
        RECT 47.800 67.900 48.200 70.200 ;
        RECT 49.400 67.900 49.800 70.200 ;
        RECT 52.400 67.900 52.800 70.200 ;
        RECT 53.400 68.900 53.800 70.200 ;
        RECT 55.000 68.900 55.400 70.200 ;
        RECT 56.900 68.000 57.300 70.200 ;
        RECT 59.800 68.300 60.200 70.200 ;
        RECT 63.800 68.900 64.200 70.200 ;
        RECT 66.200 68.300 66.600 70.200 ;
        RECT 69.500 69.900 69.900 70.200 ;
        RECT 69.400 68.200 69.900 69.900 ;
        RECT 72.500 68.200 73.000 70.200 ;
        RECT 75.800 67.900 76.200 70.200 ;
        RECT 77.400 67.900 77.800 70.200 ;
        RECT 79.000 68.900 79.400 70.200 ;
        RECT 80.600 68.900 81.000 70.200 ;
        RECT 81.400 67.900 81.800 70.200 ;
        RECT 84.600 68.900 85.000 70.200 ;
        RECT 0.600 50.800 1.000 53.100 ;
        RECT 2.200 50.800 2.600 52.100 ;
        RECT 3.800 50.800 4.200 52.100 ;
        RECT 6.200 50.800 6.600 53.100 ;
        RECT 7.000 50.800 7.400 52.100 ;
        RECT 9.100 50.800 9.500 53.100 ;
        RECT 10.200 50.800 10.600 52.100 ;
        RECT 11.800 50.800 12.200 52.100 ;
        RECT 12.600 50.800 13.000 52.100 ;
        RECT 15.800 50.800 16.200 53.100 ;
        RECT 18.200 50.800 18.600 52.700 ;
        RECT 19.800 50.800 20.200 52.100 ;
        RECT 21.900 50.800 22.300 53.100 ;
        RECT 25.400 50.800 25.800 52.700 ;
        RECT 28.600 51.100 29.100 52.800 ;
        RECT 28.700 50.800 29.100 51.100 ;
        RECT 31.700 50.800 32.200 52.800 ;
        RECT 33.400 50.800 33.800 53.100 ;
        RECT 36.400 50.800 36.800 53.100 ;
        RECT 37.400 50.800 37.800 53.100 ;
        RECT 40.600 50.800 41.000 52.100 ;
        RECT 41.400 50.800 41.800 53.100 ;
        RECT 43.800 50.800 44.200 53.100 ;
        RECT 46.200 50.800 46.600 52.100 ;
        RECT 47.800 50.800 48.200 52.100 ;
        RECT 48.600 50.800 49.000 52.100 ;
        RECT 50.200 50.800 50.600 52.100 ;
        RECT 51.000 50.800 51.400 53.100 ;
        RECT 52.600 50.800 53.000 53.100 ;
        RECT 55.000 50.800 55.400 52.100 ;
        RECT 56.600 50.800 57.000 52.100 ;
        RECT 57.400 50.800 57.800 53.100 ;
        RECT 59.000 50.800 59.400 53.100 ;
        RECT 63.000 50.800 63.400 54.100 ;
        RECT 66.400 50.800 66.800 53.100 ;
        RECT 69.400 50.800 69.800 53.100 ;
        RECT 71.000 50.800 71.400 53.100 ;
        RECT 73.400 50.800 73.800 52.700 ;
        RECT 75.300 50.800 75.700 53.100 ;
        RECT 77.400 50.800 77.800 52.100 ;
        RECT 78.200 50.800 78.600 52.100 ;
        RECT 80.300 50.800 80.700 53.100 ;
        RECT 81.400 50.800 81.800 54.100 ;
        RECT 85.400 50.800 85.800 53.100 ;
        RECT 0.200 50.200 87.800 50.800 ;
        RECT 1.400 47.900 1.800 50.200 ;
        RECT 3.000 48.900 3.400 50.200 ;
        RECT 5.100 47.900 5.500 50.200 ;
        RECT 7.800 48.300 8.200 50.200 ;
        RECT 11.000 48.300 11.400 50.200 ;
        RECT 13.700 48.000 14.100 50.200 ;
        RECT 16.600 48.300 17.000 50.200 ;
        RECT 19.000 48.900 19.400 50.200 ;
        RECT 21.100 47.900 21.500 50.200 ;
        RECT 23.000 47.900 23.400 50.200 ;
        RECT 26.200 48.300 26.600 50.200 ;
        RECT 28.600 48.900 29.000 50.200 ;
        RECT 30.200 48.900 30.600 50.200 ;
        RECT 31.800 48.300 32.200 50.200 ;
        RECT 34.200 47.900 34.600 50.200 ;
        RECT 37.200 47.900 37.600 50.200 ;
        RECT 38.200 47.900 38.600 50.200 ;
        RECT 39.800 47.900 40.200 50.200 ;
        RECT 40.600 48.900 41.000 50.200 ;
        RECT 42.200 48.900 42.600 50.200 ;
        RECT 44.600 48.300 45.000 50.200 ;
        RECT 46.200 48.900 46.600 50.200 ;
        RECT 47.800 48.900 48.200 50.200 ;
        RECT 48.600 48.900 49.000 50.200 ;
        RECT 50.200 48.900 50.600 50.200 ;
        RECT 51.000 48.900 51.400 50.200 ;
        RECT 52.600 48.900 53.000 50.200 ;
        RECT 55.000 48.300 55.400 50.200 ;
        RECT 57.400 47.900 57.800 50.200 ;
        RECT 59.800 47.900 60.200 50.200 ;
        RECT 62.200 47.900 62.600 50.200 ;
        RECT 64.600 47.900 65.000 50.200 ;
        RECT 67.600 47.900 68.000 50.200 ;
        RECT 68.600 47.900 69.000 50.200 ;
        RECT 70.200 47.900 70.600 50.200 ;
        RECT 72.600 47.900 73.000 50.200 ;
        RECT 75.800 46.900 76.200 50.200 ;
        RECT 79.000 46.900 79.400 50.200 ;
        RECT 79.800 47.900 80.200 50.200 ;
        RECT 82.200 48.900 82.600 50.200 ;
        RECT 84.300 47.900 84.700 50.200 ;
        RECT 87.000 47.900 87.400 50.200 ;
        RECT 1.400 31.100 1.900 32.800 ;
        RECT 1.500 30.800 1.900 31.100 ;
        RECT 4.500 30.800 5.000 32.800 ;
        RECT 7.800 30.800 8.200 32.700 ;
        RECT 9.400 30.800 9.800 33.100 ;
        RECT 12.600 30.800 13.000 32.700 ;
        RECT 15.000 30.800 15.400 32.100 ;
        RECT 16.600 30.800 17.000 32.100 ;
        RECT 18.200 30.800 18.600 32.700 ;
        RECT 20.900 30.800 21.300 33.100 ;
        RECT 23.000 30.800 23.400 32.100 ;
        RECT 26.200 30.800 26.600 32.100 ;
        RECT 27.000 30.800 27.400 32.100 ;
        RECT 28.600 30.800 29.000 32.100 ;
        RECT 30.200 30.800 30.600 32.100 ;
        RECT 32.600 30.800 33.000 33.100 ;
        RECT 33.400 30.800 33.800 33.100 ;
        RECT 36.400 30.800 36.800 33.100 ;
        RECT 37.700 30.800 38.100 33.100 ;
        RECT 39.800 30.800 40.200 32.100 ;
        RECT 40.600 30.800 41.000 33.100 ;
        RECT 43.800 30.800 44.200 32.700 ;
        RECT 46.500 30.800 46.900 33.100 ;
        RECT 48.600 30.800 49.000 32.100 ;
        RECT 50.200 30.800 50.600 32.100 ;
        RECT 51.300 30.800 51.700 33.100 ;
        RECT 53.400 30.800 53.800 32.100 ;
        RECT 55.800 30.800 56.200 32.700 ;
        RECT 57.400 30.800 57.800 33.100 ;
        RECT 59.800 30.800 60.200 32.700 ;
        RECT 64.600 30.800 65.000 32.700 ;
        RECT 67.000 30.800 67.400 32.100 ;
        RECT 68.600 30.800 69.000 32.100 ;
        RECT 70.200 30.800 70.600 32.700 ;
        RECT 72.600 30.800 73.000 33.100 ;
        RECT 77.400 30.800 77.800 34.100 ;
        RECT 78.200 30.800 78.600 34.100 ;
        RECT 82.200 30.800 82.600 32.700 ;
        RECT 85.400 30.800 85.800 33.100 ;
        RECT 0.200 30.200 87.800 30.800 ;
        RECT 1.500 29.900 1.900 30.200 ;
        RECT 1.400 28.200 1.900 29.900 ;
        RECT 4.500 28.200 5.000 30.200 ;
        RECT 7.800 27.900 8.200 30.200 ;
        RECT 8.600 26.900 9.000 30.200 ;
        RECT 12.600 28.300 13.000 30.200 ;
        RECT 15.000 28.900 15.400 30.200 ;
        RECT 16.600 28.900 17.000 30.200 ;
        RECT 18.200 28.300 18.600 30.200 ;
        RECT 21.400 28.300 21.800 30.200 ;
        RECT 27.000 28.300 27.400 30.200 ;
        RECT 28.600 28.900 29.000 30.200 ;
        RECT 30.200 28.900 30.600 30.200 ;
        RECT 31.800 27.900 32.200 30.200 ;
        RECT 33.400 28.300 33.800 30.200 ;
        RECT 35.800 27.900 36.200 30.200 ;
        RECT 38.800 27.900 39.200 30.200 ;
        RECT 39.800 28.900 40.200 30.200 ;
        RECT 41.400 28.900 41.800 30.200 ;
        RECT 42.500 27.900 42.900 30.200 ;
        RECT 44.600 28.900 45.000 30.200 ;
        RECT 46.200 28.300 46.600 30.200 ;
        RECT 48.900 27.900 49.300 30.200 ;
        RECT 51.000 28.900 51.400 30.200 ;
        RECT 51.800 28.900 52.200 30.200 ;
        RECT 55.800 28.300 56.200 30.200 ;
        RECT 57.400 27.900 57.800 30.200 ;
        RECT 61.400 28.900 61.800 30.200 ;
        RECT 63.000 28.900 63.400 30.200 ;
        RECT 64.600 28.300 65.000 30.200 ;
        RECT 68.600 27.900 69.000 30.200 ;
        RECT 71.000 27.900 71.400 30.200 ;
        RECT 71.800 27.900 72.200 30.200 ;
        RECT 73.400 27.900 73.800 30.200 ;
        RECT 74.200 28.900 74.600 30.200 ;
        RECT 76.100 27.900 76.500 30.200 ;
        RECT 78.200 28.900 78.600 30.200 ;
        RECT 79.000 28.900 79.400 30.200 ;
        RECT 81.400 28.300 81.800 30.200 ;
        RECT 83.800 27.900 84.200 30.200 ;
        RECT 1.400 10.800 1.800 13.100 ;
        RECT 5.400 10.800 5.800 14.100 ;
        RECT 7.000 10.800 7.400 12.700 ;
        RECT 9.400 10.800 9.800 12.100 ;
        RECT 11.500 10.800 11.900 13.100 ;
        RECT 13.400 10.800 13.800 12.700 ;
        RECT 15.800 10.800 16.200 12.100 ;
        RECT 17.400 10.800 17.800 12.100 ;
        RECT 19.000 10.800 19.400 12.700 ;
        RECT 21.400 10.800 21.800 12.100 ;
        RECT 23.000 10.800 23.400 12.100 ;
        RECT 27.000 10.800 27.400 12.700 ;
        RECT 28.900 10.800 29.300 13.100 ;
        RECT 31.000 10.800 31.400 12.100 ;
        RECT 32.600 10.800 33.000 12.700 ;
        RECT 35.800 10.800 36.200 12.100 ;
        RECT 36.600 10.800 37.000 12.100 ;
        RECT 38.200 10.800 38.600 12.100 ;
        RECT 40.600 10.800 41.000 12.700 ;
        RECT 43.300 10.800 43.700 13.000 ;
        RECT 45.400 10.800 45.800 12.100 ;
        RECT 47.000 10.800 47.400 12.100 ;
        RECT 48.600 10.800 49.000 12.700 ;
        RECT 51.800 10.800 52.200 13.100 ;
        RECT 54.800 10.800 55.200 13.100 ;
        RECT 57.400 10.800 57.800 12.700 ;
        RECT 60.300 10.800 60.700 13.000 ;
        RECT 64.600 10.800 65.000 12.700 ;
        RECT 67.200 10.800 67.600 13.100 ;
        RECT 70.200 10.800 70.600 13.100 ;
        RECT 71.000 10.800 71.400 12.100 ;
        RECT 72.600 10.800 73.000 12.900 ;
        RECT 74.500 10.800 74.900 13.100 ;
        RECT 76.600 10.800 77.000 12.100 ;
        RECT 78.200 10.800 78.600 12.700 ;
        RECT 81.700 10.800 82.100 13.000 ;
        RECT 84.600 10.800 85.000 12.100 ;
        RECT 86.200 10.800 86.600 13.100 ;
        RECT 0.200 10.200 87.800 10.800 ;
        RECT 1.400 7.900 1.800 10.200 ;
        RECT 3.900 9.900 4.300 10.200 ;
        RECT 3.800 8.200 4.300 9.900 ;
        RECT 6.900 8.200 7.400 10.200 ;
        RECT 9.400 8.300 9.800 10.200 ;
        RECT 12.900 8.000 13.300 10.200 ;
        RECT 15.900 9.900 16.300 10.200 ;
        RECT 15.800 8.200 16.300 9.900 ;
        RECT 18.900 8.200 19.400 10.200 ;
        RECT 21.400 8.200 21.900 10.200 ;
        RECT 24.500 9.900 24.900 10.200 ;
        RECT 24.500 8.200 25.000 9.900 ;
        RECT 27.800 7.900 28.200 10.200 ;
        RECT 30.200 7.900 30.600 10.200 ;
        RECT 33.100 8.000 33.500 10.200 ;
        RECT 35.800 7.900 36.200 10.200 ;
        RECT 39.000 8.300 39.400 10.200 ;
        RECT 41.400 8.900 41.800 10.200 ;
        RECT 43.800 8.300 44.200 10.200 ;
        RECT 47.000 7.900 47.400 10.200 ;
        RECT 49.400 8.300 49.800 10.200 ;
        RECT 51.000 7.900 51.400 10.200 ;
        RECT 54.200 8.900 54.600 10.200 ;
        RECT 56.600 7.900 57.000 10.200 ;
        RECT 57.400 7.900 57.800 10.200 ;
        RECT 59.000 7.900 59.400 10.200 ;
        RECT 61.400 8.900 61.800 10.200 ;
        RECT 63.000 8.900 63.400 10.200 ;
        RECT 63.800 8.900 64.200 10.200 ;
        RECT 66.200 8.300 66.600 10.200 ;
        RECT 69.500 9.900 69.900 10.200 ;
        RECT 69.400 8.200 69.900 9.900 ;
        RECT 72.500 8.200 73.000 10.200 ;
        RECT 75.100 9.900 75.500 10.200 ;
        RECT 75.000 8.200 75.500 9.900 ;
        RECT 78.100 8.200 78.600 10.200 ;
        RECT 79.800 8.900 80.200 10.200 ;
        RECT 82.200 8.300 82.600 10.200 ;
        RECT 85.400 7.900 85.800 10.200 ;
      LAYER via1 ;
        RECT 61.000 70.300 61.400 70.700 ;
        RECT 61.700 70.300 62.100 70.700 ;
        RECT 61.000 50.300 61.400 50.700 ;
        RECT 61.700 50.300 62.100 50.700 ;
        RECT 61.000 30.300 61.400 30.700 ;
        RECT 61.700 30.300 62.100 30.700 ;
        RECT 61.000 10.300 61.400 10.700 ;
        RECT 61.700 10.300 62.100 10.700 ;
      LAYER metal2 ;
        RECT 60.800 70.300 62.400 70.700 ;
        RECT 60.800 50.300 62.400 50.700 ;
        RECT 60.800 30.300 62.400 30.700 ;
        RECT 60.800 10.300 62.400 10.700 ;
      LAYER via2 ;
        RECT 61.000 70.300 61.400 70.700 ;
        RECT 61.700 70.300 62.100 70.700 ;
        RECT 61.000 50.300 61.400 50.700 ;
        RECT 61.700 50.300 62.100 50.700 ;
        RECT 61.000 30.300 61.400 30.700 ;
        RECT 61.700 30.300 62.100 30.700 ;
        RECT 61.000 10.300 61.400 10.700 ;
        RECT 61.700 10.300 62.100 10.700 ;
      LAYER metal3 ;
        RECT 60.800 70.300 62.400 70.700 ;
        RECT 60.800 50.300 62.400 50.700 ;
        RECT 60.800 30.300 62.400 30.700 ;
        RECT 60.800 10.300 62.400 10.700 ;
      LAYER via3 ;
        RECT 61.000 70.300 61.400 70.700 ;
        RECT 61.800 70.300 62.200 70.700 ;
        RECT 61.000 50.300 61.400 50.700 ;
        RECT 61.800 50.300 62.200 50.700 ;
        RECT 61.000 30.300 61.400 30.700 ;
        RECT 61.800 30.300 62.200 30.700 ;
        RECT 61.000 10.300 61.400 10.700 ;
        RECT 61.800 10.300 62.200 10.700 ;
      LAYER metal4 ;
        RECT 60.800 70.300 62.400 70.700 ;
        RECT 60.800 50.300 62.400 50.700 ;
        RECT 60.800 30.300 62.400 30.700 ;
        RECT 60.800 10.300 62.400 10.700 ;
      LAYER via4 ;
        RECT 61.000 70.300 61.400 70.700 ;
        RECT 61.700 70.300 62.100 70.700 ;
        RECT 61.000 50.300 61.400 50.700 ;
        RECT 61.700 50.300 62.100 50.700 ;
        RECT 61.000 30.300 61.400 30.700 ;
        RECT 61.700 30.300 62.100 30.700 ;
        RECT 61.000 10.300 61.400 10.700 ;
        RECT 61.700 10.300 62.100 10.700 ;
      LAYER metal5 ;
        RECT 60.800 70.200 62.400 70.700 ;
        RECT 60.800 50.200 62.400 50.700 ;
        RECT 60.800 30.200 62.400 30.700 ;
        RECT 60.800 10.200 62.400 10.700 ;
      LAYER via5 ;
        RECT 61.800 70.200 62.300 70.700 ;
        RECT 61.800 50.200 62.300 50.700 ;
        RECT 61.800 30.200 62.300 30.700 ;
        RECT 61.800 10.200 62.300 10.700 ;
      LAYER metal6 ;
        RECT 60.800 -3.000 62.400 73.000 ;
    END
  END gnd
  PIN A[0]
    PORT
      LAYER metal1 ;
        RECT 3.800 67.800 4.200 68.600 ;
        RECT 15.000 67.800 15.400 68.600 ;
        RECT 3.800 67.100 4.100 67.800 ;
        RECT 4.600 67.100 5.000 67.600 ;
        RECT 3.800 66.800 5.000 67.100 ;
        RECT 15.000 67.100 15.300 67.800 ;
        RECT 16.200 67.200 16.600 67.400 ;
        RECT 15.800 67.100 16.600 67.200 ;
        RECT 15.000 66.900 16.600 67.100 ;
        RECT 15.000 66.800 16.200 66.900 ;
        RECT 33.400 46.100 33.800 46.200 ;
        RECT 34.200 46.100 34.600 46.200 ;
        RECT 33.400 45.800 34.600 46.100 ;
        RECT 34.200 45.400 34.600 45.800 ;
      LAYER metal2 ;
        RECT 15.000 72.800 15.400 73.200 ;
        RECT 15.000 70.200 15.300 72.800 ;
        RECT 3.800 69.800 4.200 70.200 ;
        RECT 15.000 69.800 15.400 70.200 ;
        RECT 3.800 68.200 4.100 69.800 ;
        RECT 15.000 68.200 15.300 69.800 ;
        RECT 3.800 67.800 4.200 68.200 ;
        RECT 15.000 67.800 15.400 68.200 ;
        RECT 15.000 59.200 15.300 67.800 ;
        RECT 15.000 58.800 15.400 59.200 ;
        RECT 33.400 58.800 33.800 59.200 ;
        RECT 33.400 46.200 33.700 58.800 ;
        RECT 33.400 45.800 33.800 46.200 ;
      LAYER metal3 ;
        RECT 3.800 70.100 4.200 70.200 ;
        RECT 15.000 70.100 15.400 70.200 ;
        RECT 3.800 69.800 15.400 70.100 ;
        RECT 15.000 59.100 15.400 59.200 ;
        RECT 33.400 59.100 33.800 59.200 ;
        RECT 15.000 58.800 33.800 59.100 ;
    END
  END A[0]
  PIN A[1]
    PORT
      LAYER metal1 ;
        RECT 24.600 55.100 25.000 55.200 ;
        RECT 25.400 55.100 25.800 55.200 ;
        RECT 33.400 55.100 33.800 55.600 ;
        RECT 24.600 54.800 25.800 55.100 ;
        RECT 25.400 54.400 25.800 54.800 ;
        RECT 32.600 54.800 33.800 55.100 ;
        RECT 32.600 54.200 32.900 54.800 ;
        RECT 0.600 53.400 1.000 54.200 ;
        RECT 15.800 53.400 16.200 54.200 ;
        RECT 32.200 53.800 33.000 54.200 ;
        RECT 32.600 35.100 33.000 35.200 ;
        RECT 33.400 35.100 33.800 35.600 ;
        RECT 32.600 34.800 33.800 35.100 ;
      LAYER via1 ;
        RECT 0.600 53.800 1.000 54.200 ;
        RECT 15.800 53.800 16.200 54.200 ;
        RECT 32.600 53.800 33.000 54.200 ;
      LAYER metal2 ;
        RECT 0.600 54.800 1.000 55.200 ;
        RECT 24.600 54.800 25.000 55.200 ;
        RECT 0.600 54.200 0.900 54.800 ;
        RECT 0.600 53.800 1.000 54.200 ;
        RECT 15.800 53.800 16.200 54.200 ;
        RECT 0.600 52.200 0.900 53.800 ;
        RECT 15.800 52.200 16.100 53.800 ;
        RECT 24.600 52.200 24.900 54.800 ;
        RECT 32.600 53.800 33.000 54.200 ;
        RECT 32.600 52.200 32.900 53.800 ;
        RECT 0.600 51.800 1.000 52.200 ;
        RECT 15.800 51.800 16.200 52.200 ;
        RECT 24.600 51.800 25.000 52.200 ;
        RECT 32.600 51.800 33.000 52.200 ;
        RECT 32.600 35.200 32.900 51.800 ;
        RECT 32.600 34.800 33.000 35.200 ;
      LAYER metal3 ;
        RECT -2.600 55.100 -2.200 55.200 ;
        RECT 0.600 55.100 1.000 55.200 ;
        RECT -2.600 54.800 1.000 55.100 ;
        RECT 0.600 52.100 1.000 52.200 ;
        RECT 15.800 52.100 16.200 52.200 ;
        RECT 24.600 52.100 25.000 52.200 ;
        RECT 32.600 52.100 33.000 52.200 ;
        RECT 0.600 51.800 33.000 52.100 ;
    END
  END A[1]
  PIN A[2]
    PORT
      LAYER metal1 ;
        RECT 0.600 34.100 1.400 34.200 ;
        RECT 0.600 33.800 2.300 34.100 ;
        RECT 2.000 33.600 2.300 33.800 ;
        RECT 4.000 33.800 4.400 34.200 ;
        RECT 4.000 33.600 4.300 33.800 ;
        RECT 2.000 33.300 3.000 33.600 ;
        RECT 2.200 33.200 3.000 33.300 ;
        RECT 3.900 33.200 4.300 33.600 ;
        RECT 32.600 33.400 33.000 34.200 ;
        RECT 27.400 27.200 27.800 27.400 ;
        RECT 0.600 27.100 1.400 27.200 ;
        RECT 0.600 27.000 1.700 27.100 ;
        RECT 0.600 26.800 2.800 27.000 ;
        RECT 27.400 26.900 28.200 27.200 ;
        RECT 27.800 26.800 28.200 26.900 ;
        RECT 31.800 26.800 32.200 27.600 ;
        RECT 1.400 26.700 2.800 26.800 ;
        RECT 2.400 26.600 2.800 26.700 ;
        RECT 35.800 25.400 36.200 26.200 ;
      LAYER via1 ;
        RECT 32.600 33.800 33.000 34.200 ;
        RECT 35.800 25.800 36.200 26.200 ;
      LAYER metal2 ;
        RECT 0.600 33.800 1.000 34.200 ;
        RECT 32.600 33.800 33.000 34.200 ;
        RECT 0.600 27.200 0.900 33.800 ;
        RECT 2.200 33.500 2.600 33.600 ;
        RECT 3.900 33.500 4.300 33.600 ;
        RECT 2.200 33.200 4.300 33.500 ;
        RECT 32.600 28.100 32.900 33.800 ;
        RECT 31.800 27.800 32.900 28.100 ;
        RECT 31.800 27.200 32.100 27.800 ;
        RECT 0.600 26.800 1.000 27.200 ;
        RECT 27.000 27.100 27.400 27.200 ;
        RECT 27.800 27.100 28.200 27.200 ;
        RECT 27.000 26.800 28.200 27.100 ;
        RECT 31.000 27.100 31.400 27.200 ;
        RECT 31.800 27.100 32.200 27.200 ;
        RECT 31.000 26.800 32.200 27.100 ;
        RECT 35.800 26.800 36.200 27.200 ;
        RECT 35.800 26.200 36.100 26.800 ;
        RECT 35.800 25.800 36.200 26.200 ;
      LAYER metal3 ;
        RECT -2.600 27.100 -2.200 27.200 ;
        RECT 0.600 27.100 1.000 27.200 ;
        RECT 27.000 27.100 27.400 27.200 ;
        RECT 31.000 27.100 31.400 27.200 ;
        RECT 35.800 27.100 36.200 27.200 ;
        RECT -2.600 26.800 36.200 27.100 ;
    END
  END A[2]
  PIN A[3]
    PORT
      LAYER metal1 ;
        RECT 27.800 14.100 28.200 14.200 ;
        RECT 27.400 13.800 28.200 14.100 ;
        RECT 27.400 13.600 27.800 13.800 ;
        RECT 16.600 7.700 17.400 7.800 ;
        RECT 16.400 7.400 17.400 7.700 ;
        RECT 18.300 7.400 18.700 7.800 ;
        RECT 16.400 7.200 16.700 7.400 ;
        RECT 15.000 6.900 16.700 7.200 ;
        RECT 18.400 7.200 18.700 7.400 ;
        RECT 15.000 6.800 15.800 6.900 ;
        RECT 18.400 6.800 18.800 7.200 ;
        RECT 25.000 7.100 25.800 7.200 ;
        RECT 24.700 7.000 25.800 7.100 ;
        RECT 23.600 6.800 25.800 7.000 ;
        RECT 30.200 6.800 30.600 7.600 ;
        RECT 23.600 6.700 25.000 6.800 ;
        RECT 23.600 6.600 24.000 6.700 ;
        RECT 31.800 6.400 32.200 7.200 ;
      LAYER via1 ;
        RECT 27.800 13.800 28.200 14.200 ;
        RECT 16.600 7.400 17.000 7.800 ;
        RECT 25.400 6.800 25.800 7.200 ;
        RECT 31.800 6.800 32.200 7.200 ;
      LAYER metal2 ;
        RECT 27.800 13.800 28.200 14.200 ;
        RECT 27.800 8.200 28.100 13.800 ;
        RECT 18.200 7.800 18.600 8.200 ;
        RECT 25.400 7.800 25.800 8.200 ;
        RECT 27.800 7.800 28.200 8.200 ;
        RECT 30.200 7.800 30.600 8.200 ;
        RECT 31.800 7.800 32.200 8.200 ;
        RECT 16.600 7.500 18.700 7.800 ;
        RECT 16.600 7.400 17.000 7.500 ;
        RECT 18.300 7.400 18.700 7.500 ;
        RECT 25.400 7.200 25.700 7.800 ;
        RECT 30.200 7.200 30.500 7.800 ;
        RECT 31.800 7.200 32.100 7.800 ;
        RECT 25.400 6.800 25.800 7.200 ;
        RECT 30.200 6.800 30.600 7.200 ;
        RECT 31.800 6.800 32.200 7.200 ;
        RECT 30.200 -1.800 30.500 6.800 ;
        RECT 30.200 -2.200 30.600 -1.800 ;
      LAYER metal3 ;
        RECT 18.200 8.100 18.600 8.200 ;
        RECT 25.400 8.100 25.800 8.200 ;
        RECT 27.800 8.100 28.200 8.200 ;
        RECT 30.200 8.100 30.600 8.200 ;
        RECT 31.800 8.100 32.200 8.200 ;
        RECT 18.200 7.800 32.200 8.100 ;
    END
  END A[3]
  PIN A[4]
    PORT
      LAYER metal1 ;
        RECT 56.600 7.100 57.000 7.600 ;
        RECT 57.400 7.100 57.800 7.600 ;
        RECT 56.600 6.800 57.800 7.100 ;
      LAYER via1 ;
        RECT 57.400 6.800 57.800 7.200 ;
      LAYER metal2 ;
        RECT 57.400 6.800 57.800 7.200 ;
        RECT 57.400 -1.800 57.700 6.800 ;
        RECT 57.400 -2.200 57.800 -1.800 ;
    END
  END A[4]
  PIN A[5]
    PORT
      LAYER metal1 ;
        RECT 67.000 47.100 67.400 47.200 ;
        RECT 68.600 47.100 69.000 47.200 ;
        RECT 67.000 46.800 69.000 47.100 ;
        RECT 67.000 46.400 67.400 46.800 ;
        RECT 83.800 26.800 84.200 27.600 ;
        RECT 86.200 13.400 86.600 14.200 ;
      LAYER via1 ;
        RECT 68.600 46.800 69.000 47.200 ;
        RECT 86.200 13.800 86.600 14.200 ;
      LAYER metal2 ;
        RECT 68.600 46.800 69.000 47.200 ;
        RECT 68.600 39.200 68.900 46.800 ;
        RECT 68.600 38.800 69.000 39.200 ;
        RECT 83.000 38.800 83.400 39.200 ;
        RECT 83.000 35.100 83.300 38.800 ;
        RECT 83.000 34.800 84.100 35.100 ;
        RECT 83.800 27.200 84.100 34.800 ;
        RECT 83.800 26.800 84.200 27.200 ;
        RECT 83.800 20.200 84.100 26.800 ;
        RECT 83.800 19.800 84.200 20.200 ;
        RECT 86.200 19.800 86.600 20.200 ;
        RECT 86.200 15.200 86.500 19.800 ;
        RECT 86.200 14.800 86.600 15.200 ;
        RECT 86.200 14.200 86.500 14.800 ;
        RECT 86.200 13.800 86.600 14.200 ;
      LAYER metal3 ;
        RECT 68.600 39.100 69.000 39.200 ;
        RECT 83.000 39.100 83.400 39.200 ;
        RECT 68.600 38.800 83.400 39.100 ;
        RECT 83.800 20.100 84.200 20.200 ;
        RECT 86.200 20.100 86.600 20.200 ;
        RECT 83.800 19.800 86.600 20.100 ;
        RECT 86.200 15.100 86.600 15.200 ;
        RECT 90.200 15.100 90.600 15.200 ;
        RECT 86.200 14.800 90.600 15.100 ;
    END
  END A[5]
  PIN A[6]
    PORT
      LAYER metal1 ;
        RECT 51.000 53.400 51.400 54.200 ;
        RECT 55.400 47.200 55.800 47.400 ;
        RECT 55.400 46.900 56.200 47.200 ;
        RECT 55.800 46.800 56.200 46.900 ;
        RECT 59.800 47.100 60.200 47.600 ;
        RECT 62.200 47.100 62.600 47.600 ;
        RECT 59.800 46.800 62.600 47.100 ;
        RECT 59.800 46.200 60.100 46.800 ;
        RECT 59.800 45.800 60.200 46.200 ;
      LAYER via1 ;
        RECT 51.000 53.800 51.400 54.200 ;
      LAYER metal2 ;
        RECT 51.000 73.100 51.400 73.200 ;
        RECT 51.000 72.800 52.100 73.100 ;
        RECT 51.800 54.200 52.100 72.800 ;
        RECT 51.000 54.100 51.400 54.200 ;
        RECT 51.800 54.100 52.200 54.200 ;
        RECT 51.000 53.800 52.200 54.100 ;
        RECT 55.800 53.800 56.200 54.200 ;
        RECT 55.800 47.200 56.100 53.800 ;
        RECT 55.800 47.100 56.200 47.200 ;
        RECT 56.600 47.100 57.000 47.200 ;
        RECT 55.800 46.800 57.000 47.100 ;
        RECT 59.800 46.800 60.200 47.200 ;
        RECT 59.800 46.200 60.100 46.800 ;
        RECT 59.800 45.800 60.200 46.200 ;
      LAYER via2 ;
        RECT 51.800 53.800 52.200 54.200 ;
        RECT 56.600 46.800 57.000 47.200 ;
      LAYER metal3 ;
        RECT 51.800 54.100 52.200 54.200 ;
        RECT 55.800 54.100 56.200 54.200 ;
        RECT 51.800 53.800 56.200 54.100 ;
        RECT 56.600 47.100 57.000 47.200 ;
        RECT 59.800 47.100 60.200 47.200 ;
        RECT 56.600 46.800 60.200 47.100 ;
    END
  END A[6]
  PIN A[7]
    PORT
      LAYER metal1 ;
        RECT 63.000 68.100 63.400 68.200 ;
        RECT 63.800 68.100 64.200 68.600 ;
        RECT 63.000 67.800 64.200 68.100 ;
        RECT 70.200 67.700 71.000 67.800 ;
        RECT 70.000 67.400 71.000 67.700 ;
        RECT 71.900 67.400 72.300 67.800 ;
        RECT 59.400 67.200 59.800 67.400 ;
        RECT 70.000 67.200 70.300 67.400 ;
        RECT 58.200 67.100 58.600 67.200 ;
        RECT 59.000 67.100 59.800 67.200 ;
        RECT 58.200 66.900 59.800 67.100 ;
        RECT 68.600 66.900 70.300 67.200 ;
        RECT 72.000 67.200 72.300 67.400 ;
        RECT 58.200 66.800 59.400 66.900 ;
        RECT 68.600 66.800 69.400 66.900 ;
        RECT 72.000 66.800 72.400 67.200 ;
        RECT 58.200 66.400 58.600 66.800 ;
        RECT 64.600 45.400 65.000 46.200 ;
      LAYER via1 ;
        RECT 70.200 67.400 70.600 67.800 ;
        RECT 59.000 66.800 59.400 67.200 ;
        RECT 64.600 45.800 65.000 46.200 ;
      LAYER metal2 ;
        RECT 63.000 72.800 63.400 73.200 ;
        RECT 63.000 68.200 63.300 72.800 ;
        RECT 63.000 67.800 63.400 68.200 ;
        RECT 63.000 67.200 63.300 67.800 ;
        RECT 70.200 67.500 72.300 67.800 ;
        RECT 70.200 67.400 70.600 67.500 ;
        RECT 71.900 67.400 72.300 67.500 ;
        RECT 58.200 67.100 58.600 67.200 ;
        RECT 59.000 67.100 59.400 67.200 ;
        RECT 58.200 66.800 59.400 67.100 ;
        RECT 63.000 66.800 63.400 67.200 ;
        RECT 67.800 67.100 68.200 67.200 ;
        RECT 68.600 67.100 69.000 67.200 ;
        RECT 67.800 66.800 69.000 67.100 ;
        RECT 64.600 46.800 65.000 47.200 ;
        RECT 64.600 46.200 64.900 46.800 ;
        RECT 64.600 45.800 65.000 46.200 ;
      LAYER metal3 ;
        RECT 58.200 67.100 58.600 67.200 ;
        RECT 63.000 67.100 63.400 67.200 ;
        RECT 64.600 67.100 65.000 67.200 ;
        RECT 67.800 67.100 68.200 67.200 ;
        RECT 58.200 66.800 68.200 67.100 ;
        RECT 64.600 47.800 65.000 48.200 ;
        RECT 64.600 47.200 64.900 47.800 ;
        RECT 64.600 46.800 65.000 47.200 ;
      LAYER via3 ;
        RECT 64.600 66.800 65.000 67.200 ;
      LAYER metal4 ;
        RECT 64.600 66.800 65.000 67.200 ;
        RECT 64.600 48.200 64.900 66.800 ;
        RECT 64.600 47.800 65.000 48.200 ;
    END
  END A[7]
  PIN B[0]
    PORT
      LAYER metal1 ;
        RECT 8.600 67.800 9.000 68.600 ;
        RECT 0.600 66.800 1.000 67.600 ;
        RECT 16.600 65.800 17.000 66.600 ;
        RECT 6.200 64.400 6.600 65.200 ;
      LAYER via1 ;
        RECT 6.200 64.800 6.600 65.200 ;
      LAYER metal2 ;
        RECT 8.600 67.800 9.000 68.200 ;
        RECT 0.600 66.800 1.000 67.200 ;
        RECT 0.600 65.200 0.900 66.800 ;
        RECT 8.600 65.200 8.900 67.800 ;
        RECT 16.600 65.800 17.000 66.200 ;
        RECT 16.600 65.200 16.900 65.800 ;
        RECT 0.600 64.800 1.000 65.200 ;
        RECT 5.400 65.100 5.800 65.200 ;
        RECT 6.200 65.100 6.600 65.200 ;
        RECT 5.400 64.800 6.600 65.100 ;
        RECT 8.600 64.800 9.000 65.200 ;
        RECT 16.600 64.800 17.000 65.200 ;
      LAYER metal3 ;
        RECT -2.600 65.100 -2.200 65.200 ;
        RECT 0.600 65.100 1.000 65.200 ;
        RECT 5.400 65.100 5.800 65.200 ;
        RECT 8.600 65.100 9.000 65.200 ;
        RECT 16.600 65.100 17.000 65.200 ;
        RECT -2.600 64.800 17.000 65.100 ;
    END
  END B[0]
  PIN B[1]
    PORT
      LAYER metal1 ;
        RECT 29.600 54.300 30.000 54.400 ;
        RECT 28.600 54.200 30.000 54.300 ;
        RECT 2.200 53.800 2.600 54.200 ;
        RECT 2.200 53.200 2.500 53.800 ;
        RECT 6.200 53.400 6.600 54.200 ;
        RECT 23.800 54.100 24.200 54.200 ;
        RECT 24.600 54.100 25.000 54.200 ;
        RECT 23.800 53.800 25.400 54.100 ;
        RECT 27.800 54.000 30.000 54.200 ;
        RECT 27.800 53.900 28.900 54.000 ;
        RECT 27.800 53.800 28.600 53.900 ;
        RECT 25.000 53.600 25.400 53.800 ;
        RECT 2.200 52.400 2.600 53.200 ;
        RECT 12.600 52.400 13.000 53.200 ;
      LAYER via1 ;
        RECT 6.200 53.800 6.600 54.200 ;
        RECT 12.600 52.800 13.000 53.200 ;
      LAYER metal2 ;
        RECT 27.800 54.800 28.200 55.200 ;
        RECT 27.800 54.200 28.100 54.800 ;
        RECT 2.200 53.800 2.600 54.200 ;
        RECT 6.200 53.800 6.600 54.200 ;
        RECT 23.800 53.800 24.200 54.200 ;
        RECT 27.800 53.800 28.200 54.200 ;
        RECT 2.200 53.200 2.500 53.800 ;
        RECT 6.200 53.200 6.500 53.800 ;
        RECT 23.800 53.200 24.100 53.800 ;
        RECT 2.200 52.800 2.600 53.200 ;
        RECT 6.200 52.800 6.600 53.200 ;
        RECT 11.800 53.100 12.200 53.200 ;
        RECT 12.600 53.100 13.000 53.200 ;
        RECT 11.800 52.800 13.000 53.100 ;
        RECT 23.800 52.800 24.200 53.200 ;
      LAYER metal3 ;
        RECT 27.800 54.800 28.200 55.200 ;
        RECT 23.800 54.100 24.200 54.200 ;
        RECT 27.800 54.100 28.100 54.800 ;
        RECT 23.800 53.800 28.100 54.100 ;
        RECT -2.600 53.100 -2.200 53.200 ;
        RECT 2.200 53.100 2.600 53.200 ;
        RECT 6.200 53.100 6.600 53.200 ;
        RECT 11.800 53.100 12.200 53.200 ;
        RECT 23.800 53.100 24.200 53.200 ;
        RECT -2.600 52.800 24.200 53.100 ;
    END
  END B[1]
  PIN B[2]
    PORT
      LAYER metal1 ;
        RECT 5.000 33.800 5.800 34.200 ;
        RECT 27.000 32.400 27.400 33.200 ;
        RECT 28.600 27.800 29.000 28.600 ;
        RECT 5.000 26.800 5.800 27.200 ;
        RECT 27.000 26.100 27.400 26.600 ;
        RECT 28.600 26.100 29.000 26.200 ;
        RECT 27.000 25.800 29.000 26.100 ;
      LAYER via1 ;
        RECT 5.400 33.800 5.800 34.200 ;
        RECT 27.000 32.800 27.400 33.200 ;
        RECT 5.400 26.800 5.800 27.200 ;
        RECT 28.600 25.800 29.000 26.200 ;
      LAYER metal2 ;
        RECT 5.400 33.800 5.800 34.200 ;
        RECT 5.400 30.200 5.700 33.800 ;
        RECT 27.000 32.800 27.400 33.200 ;
        RECT 27.000 30.200 27.300 32.800 ;
        RECT 5.400 29.800 5.800 30.200 ;
        RECT 27.000 29.800 27.400 30.200 ;
        RECT 28.600 29.800 29.000 30.200 ;
        RECT 5.400 29.200 5.700 29.800 ;
        RECT 5.400 28.800 5.800 29.200 ;
        RECT 5.400 27.200 5.700 28.800 ;
        RECT 28.600 28.200 28.900 29.800 ;
        RECT 28.600 27.800 29.000 28.200 ;
        RECT 5.400 26.800 5.800 27.200 ;
        RECT 28.600 26.200 28.900 27.800 ;
        RECT 28.600 25.800 29.000 26.200 ;
      LAYER metal3 ;
        RECT 5.400 30.100 5.800 30.200 ;
        RECT 27.000 30.100 27.400 30.200 ;
        RECT 28.600 30.100 29.000 30.200 ;
        RECT 5.400 29.800 29.000 30.100 ;
        RECT -2.600 29.100 -2.200 29.200 ;
        RECT 5.400 29.100 5.800 29.200 ;
        RECT -2.600 28.800 5.800 29.100 ;
    END
  END B[2]
  PIN B[3]
    PORT
      LAYER metal1 ;
        RECT 27.000 14.400 27.400 15.200 ;
        RECT 36.600 12.400 37.000 13.200 ;
        RECT 19.400 7.100 20.200 7.200 ;
        RECT 20.600 7.100 21.400 7.200 ;
        RECT 19.400 6.800 21.400 7.100 ;
        RECT 27.800 6.800 28.200 7.600 ;
        RECT 32.800 6.900 33.200 7.000 ;
        RECT 20.600 6.200 20.900 6.800 ;
        RECT 32.700 6.600 33.200 6.900 ;
        RECT 32.700 6.200 33.000 6.600 ;
        RECT 20.600 5.800 21.000 6.200 ;
        RECT 32.600 5.800 33.000 6.200 ;
      LAYER via1 ;
        RECT 27.000 14.800 27.400 15.200 ;
        RECT 36.600 12.800 37.000 13.200 ;
      LAYER metal2 ;
        RECT 27.000 14.800 27.400 15.200 ;
        RECT 27.000 7.200 27.300 14.800 ;
        RECT 36.600 12.800 37.000 13.200 ;
        RECT 36.600 7.200 36.900 12.800 ;
        RECT 20.600 6.800 21.000 7.200 ;
        RECT 27.000 7.100 27.400 7.200 ;
        RECT 27.800 7.100 28.200 7.200 ;
        RECT 27.000 6.800 28.200 7.100 ;
        RECT 32.600 6.800 33.000 7.200 ;
        RECT 36.600 6.800 37.000 7.200 ;
        RECT 20.600 6.200 20.900 6.800 ;
        RECT 32.600 6.200 32.900 6.800 ;
        RECT 20.600 5.800 21.000 6.200 ;
        RECT 32.600 5.800 33.000 6.200 ;
        RECT 32.600 -1.800 32.900 5.800 ;
        RECT 32.600 -2.200 33.000 -1.800 ;
      LAYER metal3 ;
        RECT 20.600 7.100 21.000 7.200 ;
        RECT 27.000 7.100 27.400 7.200 ;
        RECT 32.600 7.100 33.000 7.200 ;
        RECT 36.600 7.100 37.000 7.200 ;
        RECT 20.600 6.800 37.000 7.100 ;
    END
  END B[3]
  PIN B[4]
    PORT
      LAYER metal1 ;
        RECT 54.200 7.800 54.600 8.600 ;
        RECT 59.800 8.100 60.200 8.200 ;
        RECT 61.400 8.100 61.800 8.600 ;
        RECT 59.800 7.800 61.800 8.100 ;
        RECT 54.200 5.100 54.600 5.200 ;
        RECT 55.000 5.100 55.400 5.200 ;
        RECT 54.200 4.800 55.400 5.100 ;
        RECT 55.000 3.800 55.400 4.800 ;
      LAYER metal2 ;
        RECT 54.200 7.800 54.600 8.200 ;
        RECT 59.800 7.800 60.200 8.200 ;
        RECT 54.200 7.200 54.500 7.800 ;
        RECT 59.800 7.200 60.100 7.800 ;
        RECT 54.200 6.800 54.600 7.200 ;
        RECT 59.800 6.800 60.200 7.200 ;
        RECT 54.200 5.200 54.500 6.800 ;
        RECT 54.200 4.800 54.600 5.200 ;
        RECT 55.000 3.800 55.400 4.200 ;
        RECT 55.000 -1.800 55.300 3.800 ;
        RECT 55.000 -2.200 55.400 -1.800 ;
      LAYER metal3 ;
        RECT 54.200 7.100 54.600 7.200 ;
        RECT 59.800 7.100 60.200 7.200 ;
        RECT 54.200 6.800 60.200 7.100 ;
    END
  END B[4]
  PIN B[5]
    PORT
      LAYER metal1 ;
        RECT 79.000 67.800 79.400 68.600 ;
        RECT 84.600 67.800 85.000 68.600 ;
        RECT 85.400 25.100 85.800 25.200 ;
        RECT 86.200 25.100 86.600 25.200 ;
        RECT 85.400 24.800 86.600 25.100 ;
        RECT 85.400 24.400 85.800 24.800 ;
      LAYER via1 ;
        RECT 86.200 24.800 86.600 25.200 ;
      LAYER metal2 ;
        RECT 79.000 68.100 79.400 68.200 ;
        RECT 79.800 68.100 80.200 68.200 ;
        RECT 79.000 67.800 80.200 68.100 ;
        RECT 84.600 67.800 85.000 68.200 ;
        RECT 84.600 56.200 84.900 67.800 ;
        RECT 84.600 55.800 85.000 56.200 ;
        RECT 86.200 41.800 86.600 42.200 ;
        RECT 86.200 25.200 86.500 41.800 ;
        RECT 86.200 24.800 86.600 25.200 ;
      LAYER via2 ;
        RECT 79.800 67.800 80.200 68.200 ;
      LAYER metal3 ;
        RECT 79.800 68.100 80.200 68.200 ;
        RECT 84.600 68.100 85.000 68.200 ;
        RECT 79.800 67.800 85.000 68.100 ;
        RECT 84.600 56.100 85.000 56.200 ;
        RECT 87.000 56.100 87.400 56.200 ;
        RECT 90.200 56.100 90.600 56.200 ;
        RECT 84.600 55.800 90.600 56.100 ;
        RECT 86.200 42.100 86.600 42.200 ;
        RECT 87.000 42.100 87.400 42.200 ;
        RECT 86.200 41.800 87.400 42.100 ;
      LAYER via3 ;
        RECT 87.000 55.800 87.400 56.200 ;
        RECT 87.000 41.800 87.400 42.200 ;
      LAYER metal4 ;
        RECT 87.000 55.800 87.400 56.200 ;
        RECT 87.000 42.200 87.300 55.800 ;
        RECT 87.000 41.800 87.400 42.200 ;
    END
  END B[5]
  PIN B[6]
    PORT
      LAYER metal1 ;
        RECT 52.600 53.400 53.000 54.200 ;
        RECT 56.600 53.800 57.000 54.200 ;
        RECT 56.600 53.200 56.900 53.800 ;
        RECT 56.600 52.400 57.000 53.200 ;
        RECT 55.000 45.800 55.400 46.600 ;
        RECT 58.200 44.400 58.600 45.200 ;
      LAYER via1 ;
        RECT 52.600 53.800 53.000 54.200 ;
        RECT 58.200 44.800 58.600 45.200 ;
      LAYER metal2 ;
        RECT 53.400 72.800 53.800 73.200 ;
        RECT 53.400 70.200 53.700 72.800 ;
        RECT 53.400 69.800 53.800 70.200 ;
        RECT 56.600 69.800 57.000 70.200 ;
        RECT 56.600 54.200 56.900 69.800 ;
        RECT 52.600 53.800 53.000 54.200 ;
        RECT 56.600 53.800 57.000 54.200 ;
        RECT 52.600 53.200 52.900 53.800 ;
        RECT 56.600 53.200 56.900 53.800 ;
        RECT 52.600 52.800 53.000 53.200 ;
        RECT 55.000 52.800 55.400 53.200 ;
        RECT 56.600 52.800 57.000 53.200 ;
        RECT 58.200 52.800 58.600 53.200 ;
        RECT 55.000 46.200 55.300 52.800 ;
        RECT 55.000 45.800 55.400 46.200 ;
        RECT 58.200 45.200 58.500 52.800 ;
        RECT 58.200 44.800 58.600 45.200 ;
      LAYER metal3 ;
        RECT 53.400 70.100 53.800 70.200 ;
        RECT 56.600 70.100 57.000 70.200 ;
        RECT 53.400 69.800 57.000 70.100 ;
        RECT 52.600 53.100 53.000 53.200 ;
        RECT 55.000 53.100 55.400 53.200 ;
        RECT 56.600 53.100 57.000 53.200 ;
        RECT 58.200 53.100 58.600 53.200 ;
        RECT 52.600 52.800 58.600 53.100 ;
    END
  END B[6]
  PIN B[7]
    PORT
      LAYER metal1 ;
        RECT 57.200 66.900 57.600 67.000 ;
        RECT 57.200 66.600 57.700 66.900 ;
        RECT 73.000 66.800 73.800 67.200 ;
        RECT 57.400 66.200 57.700 66.600 ;
        RECT 57.400 65.800 57.800 66.200 ;
        RECT 59.000 66.100 59.400 66.200 ;
        RECT 59.800 66.100 60.200 66.600 ;
        RECT 59.000 65.800 60.200 66.100 ;
        RECT 66.200 65.800 66.600 66.600 ;
      LAYER via1 ;
        RECT 73.400 66.800 73.800 67.200 ;
      LAYER metal2 ;
        RECT 71.000 72.800 71.400 73.200 ;
        RECT 71.000 70.200 71.300 72.800 ;
        RECT 71.000 69.800 71.400 70.200 ;
        RECT 73.400 69.800 73.800 70.200 ;
        RECT 73.400 67.200 73.700 69.800 ;
        RECT 73.400 66.800 73.800 67.200 ;
        RECT 73.400 66.200 73.700 66.800 ;
        RECT 57.400 66.100 57.800 66.200 ;
        RECT 58.200 66.100 58.600 66.200 ;
        RECT 57.400 65.800 58.600 66.100 ;
        RECT 59.000 66.100 59.400 66.200 ;
        RECT 59.800 66.100 60.200 66.200 ;
        RECT 59.000 65.800 60.200 66.100 ;
        RECT 65.400 66.100 65.800 66.200 ;
        RECT 66.200 66.100 66.600 66.200 ;
        RECT 65.400 65.800 66.600 66.100 ;
        RECT 73.400 65.800 73.800 66.200 ;
      LAYER via2 ;
        RECT 58.200 65.800 58.600 66.200 ;
        RECT 59.800 65.800 60.200 66.200 ;
      LAYER metal3 ;
        RECT 71.000 70.100 71.400 70.200 ;
        RECT 73.400 70.100 73.800 70.200 ;
        RECT 71.000 69.800 73.800 70.100 ;
        RECT 58.200 66.100 58.600 66.200 ;
        RECT 59.800 66.100 60.200 66.200 ;
        RECT 65.400 66.100 65.800 66.200 ;
        RECT 73.400 66.100 73.800 66.200 ;
        RECT 58.200 65.800 73.800 66.100 ;
    END
  END B[7]
  PIN ALU_Sel[0]
    PORT
      LAYER metal1 ;
        RECT 29.400 66.800 29.800 67.600 ;
        RECT 35.800 66.100 36.200 66.200 ;
        RECT 36.600 66.100 37.000 66.600 ;
        RECT 35.800 65.800 37.000 66.100 ;
        RECT 43.800 53.400 44.200 54.200 ;
        RECT 40.600 52.400 41.000 53.200 ;
      LAYER via1 ;
        RECT 43.800 53.800 44.200 54.200 ;
        RECT 40.600 52.800 41.000 53.200 ;
      LAYER metal2 ;
        RECT 30.200 72.800 30.600 73.200 ;
        RECT 30.200 69.200 30.500 72.800 ;
        RECT 30.200 69.100 30.600 69.200 ;
        RECT 29.400 68.800 30.600 69.100 ;
        RECT 35.800 68.800 36.200 69.200 ;
        RECT 40.600 68.800 41.000 69.200 ;
        RECT 29.400 67.200 29.700 68.800 ;
        RECT 29.400 66.800 29.800 67.200 ;
        RECT 35.800 66.200 36.100 68.800 ;
        RECT 35.800 65.800 36.200 66.200 ;
        RECT 40.600 54.200 40.900 68.800 ;
        RECT 40.600 53.800 41.000 54.200 ;
        RECT 43.000 54.100 43.400 54.200 ;
        RECT 43.800 54.100 44.200 54.200 ;
        RECT 43.000 53.800 44.200 54.100 ;
        RECT 40.600 53.200 40.900 53.800 ;
        RECT 40.600 52.800 41.000 53.200 ;
      LAYER via2 ;
        RECT 30.200 68.800 30.600 69.200 ;
      LAYER metal3 ;
        RECT 30.200 69.100 30.600 69.200 ;
        RECT 35.800 69.100 36.200 69.200 ;
        RECT 40.600 69.100 41.000 69.200 ;
        RECT 30.200 68.800 41.000 69.100 ;
        RECT 40.600 54.100 41.000 54.200 ;
        RECT 43.000 54.100 43.400 54.200 ;
        RECT 40.600 53.800 43.400 54.100 ;
    END
  END ALU_Sel[0]
  PIN ALU_Sel[1]
    PORT
      LAYER metal1 ;
        RECT 34.200 66.800 34.600 67.600 ;
        RECT 31.000 64.400 31.400 65.200 ;
        RECT 37.400 53.400 37.800 54.200 ;
      LAYER via1 ;
        RECT 31.000 64.800 31.400 65.200 ;
        RECT 37.400 53.800 37.800 54.200 ;
      LAYER metal2 ;
        RECT 32.600 72.800 33.000 73.200 ;
        RECT 32.600 70.200 32.900 72.800 ;
        RECT 32.600 69.800 33.000 70.200 ;
        RECT 34.200 69.800 34.600 70.200 ;
        RECT 34.200 67.200 34.500 69.800 ;
        RECT 34.200 66.800 34.600 67.200 ;
        RECT 31.000 64.800 31.400 65.200 ;
        RECT 31.000 64.200 31.300 64.800 ;
        RECT 34.200 64.200 34.500 66.800 ;
        RECT 31.000 63.800 31.400 64.200 ;
        RECT 34.200 63.800 34.600 64.200 ;
        RECT 37.400 63.800 37.800 64.200 ;
        RECT 37.400 54.200 37.700 63.800 ;
        RECT 37.400 53.800 37.800 54.200 ;
      LAYER metal3 ;
        RECT 32.600 70.100 33.000 70.200 ;
        RECT 34.200 70.100 34.600 70.200 ;
        RECT 32.600 69.800 34.600 70.100 ;
        RECT 31.000 64.100 31.400 64.200 ;
        RECT 34.200 64.100 34.600 64.200 ;
        RECT 37.400 64.100 37.800 64.200 ;
        RECT 31.000 63.800 37.800 64.100 ;
    END
  END ALU_Sel[1]
  PIN ALU_Sel[2]
    PORT
      LAYER metal1 ;
        RECT 22.200 67.800 22.600 68.600 ;
        RECT 21.000 67.200 21.400 67.400 ;
        RECT 21.000 67.100 21.800 67.200 ;
        RECT 22.200 67.100 22.600 67.200 ;
        RECT 21.000 66.900 22.600 67.100 ;
        RECT 21.400 66.800 22.600 66.900 ;
        RECT 42.200 66.800 42.600 67.600 ;
        RECT 46.200 52.400 46.600 53.200 ;
        RECT 40.600 47.800 41.000 48.600 ;
        RECT 46.200 47.800 46.600 48.600 ;
        RECT 44.600 46.100 45.000 46.600 ;
        RECT 46.200 46.100 46.600 46.200 ;
        RECT 44.600 45.800 46.600 46.100 ;
      LAYER via1 ;
        RECT 22.200 66.800 22.600 67.200 ;
        RECT 46.200 52.800 46.600 53.200 ;
        RECT 46.200 45.800 46.600 46.200 ;
      LAYER metal2 ;
        RECT 22.200 72.800 22.600 73.200 ;
        RECT 22.200 68.200 22.500 72.800 ;
        RECT 22.200 67.800 22.600 68.200 ;
        RECT 22.200 67.200 22.500 67.800 ;
        RECT 22.200 66.800 22.600 67.200 ;
        RECT 42.200 66.800 42.600 67.200 ;
        RECT 22.200 63.200 22.500 66.800 ;
        RECT 42.200 64.100 42.500 66.800 ;
        RECT 41.400 63.800 42.500 64.100 ;
        RECT 41.400 63.200 41.700 63.800 ;
        RECT 22.200 62.800 22.600 63.200 ;
        RECT 41.400 62.800 41.800 63.200 ;
        RECT 41.400 48.200 41.700 62.800 ;
        RECT 46.200 52.800 46.600 53.200 ;
        RECT 46.200 48.200 46.500 52.800 ;
        RECT 40.600 48.100 41.000 48.200 ;
        RECT 41.400 48.100 41.800 48.200 ;
        RECT 40.600 47.800 41.800 48.100 ;
        RECT 46.200 47.800 46.600 48.200 ;
        RECT 46.200 46.200 46.500 47.800 ;
        RECT 46.200 45.800 46.600 46.200 ;
      LAYER via2 ;
        RECT 41.400 47.800 41.800 48.200 ;
      LAYER metal3 ;
        RECT 22.200 63.100 22.600 63.200 ;
        RECT 41.400 63.100 41.800 63.200 ;
        RECT 22.200 62.800 41.800 63.100 ;
        RECT 41.400 48.100 41.800 48.200 ;
        RECT 46.200 48.100 46.600 48.200 ;
        RECT 41.400 47.800 46.600 48.100 ;
    END
  END ALU_Sel[2]
  PIN ALU_Out[0]
    PORT
      LAYER metal1 ;
        RECT 48.600 66.200 49.000 69.900 ;
        RECT 48.700 65.100 49.000 66.200 ;
        RECT 48.600 61.100 49.000 65.100 ;
      LAYER via1 ;
        RECT 48.600 68.800 49.000 69.200 ;
      LAYER metal2 ;
        RECT 47.800 73.100 48.200 73.200 ;
        RECT 47.800 72.800 48.900 73.100 ;
        RECT 48.600 69.200 48.900 72.800 ;
        RECT 48.600 68.800 49.000 69.200 ;
    END
  END ALU_Out[0]
  PIN ALU_Out[1]
    PORT
      LAYER metal1 ;
        RECT 0.600 46.200 1.000 49.900 ;
        RECT 0.600 45.100 0.900 46.200 ;
        RECT 0.600 41.100 1.000 45.100 ;
      LAYER via1 ;
        RECT 0.600 43.800 1.000 44.200 ;
      LAYER metal2 ;
        RECT 0.600 44.800 1.000 45.200 ;
        RECT 0.600 44.200 0.900 44.800 ;
        RECT 0.600 43.800 1.000 44.200 ;
      LAYER metal3 ;
        RECT -2.600 45.100 -2.200 45.200 ;
        RECT 0.600 45.100 1.000 45.200 ;
        RECT -2.600 44.800 1.000 45.100 ;
    END
  END ALU_Out[1]
  PIN ALU_Out[2]
    PORT
      LAYER metal1 ;
        RECT 0.600 15.900 1.000 19.900 ;
        RECT 0.600 14.800 0.900 15.900 ;
        RECT 0.600 11.100 1.000 14.800 ;
      LAYER via1 ;
        RECT 0.600 13.800 1.000 14.200 ;
      LAYER metal2 ;
        RECT 0.600 14.800 1.000 15.200 ;
        RECT 0.600 14.200 0.900 14.800 ;
        RECT 0.600 13.800 1.000 14.200 ;
      LAYER metal3 ;
        RECT -2.600 15.100 -2.200 15.200 ;
        RECT 0.600 15.100 1.000 15.200 ;
        RECT -2.600 14.800 1.000 15.100 ;
    END
  END ALU_Out[2]
  PIN ALU_Out[3]
    PORT
      LAYER metal1 ;
        RECT 0.600 6.200 1.000 9.900 ;
        RECT 0.600 5.100 0.900 6.200 ;
        RECT 0.600 1.100 1.000 5.100 ;
      LAYER via1 ;
        RECT 0.600 3.800 1.000 4.200 ;
      LAYER metal2 ;
        RECT 0.600 4.800 1.000 5.200 ;
        RECT 0.600 4.200 0.900 4.800 ;
        RECT 0.600 3.800 1.000 4.200 ;
      LAYER metal3 ;
        RECT -2.600 5.100 -2.200 5.200 ;
        RECT 0.600 5.100 1.000 5.200 ;
        RECT -2.600 4.800 1.000 5.100 ;
    END
  END ALU_Out[3]
  PIN ALU_Out[4]
    PORT
      LAYER metal1 ;
        RECT 35.000 6.200 35.400 9.900 ;
        RECT 35.000 5.100 35.300 6.200 ;
        RECT 35.000 1.100 35.400 5.100 ;
      LAYER via1 ;
        RECT 35.000 1.800 35.400 2.200 ;
      LAYER metal2 ;
        RECT 35.000 1.800 35.400 2.200 ;
        RECT 35.000 -1.900 35.300 1.800 ;
        RECT 35.800 -1.900 36.200 -1.800 ;
        RECT 35.000 -2.200 36.200 -1.900 ;
    END
  END ALU_Out[4]
  PIN ALU_Out[5]
    PORT
      LAYER metal1 ;
        RECT 86.200 6.200 86.600 9.900 ;
        RECT 86.300 5.100 86.600 6.200 ;
        RECT 86.200 1.100 86.600 5.100 ;
      LAYER via1 ;
        RECT 86.200 1.800 86.600 2.200 ;
      LAYER metal2 ;
        RECT 86.200 1.800 86.600 2.200 ;
        RECT 85.400 -1.900 85.800 -1.800 ;
        RECT 86.200 -1.900 86.500 1.800 ;
        RECT 85.400 -2.200 86.500 -1.900 ;
    END
  END ALU_Out[5]
  PIN ALU_Out[6]
    PORT
      LAYER metal1 ;
        RECT 86.200 35.900 86.600 39.900 ;
        RECT 86.300 34.800 86.600 35.900 ;
        RECT 86.200 34.100 86.600 34.800 ;
        RECT 87.000 34.100 87.400 34.200 ;
        RECT 86.200 33.800 87.400 34.100 ;
        RECT 86.200 31.100 86.600 33.800 ;
      LAYER via1 ;
        RECT 87.000 33.800 87.400 34.200 ;
      LAYER metal2 ;
        RECT 87.000 34.800 87.400 35.200 ;
        RECT 87.000 34.200 87.300 34.800 ;
        RECT 87.000 33.800 87.400 34.200 ;
      LAYER metal3 ;
        RECT 87.000 35.100 87.400 35.200 ;
        RECT 90.200 35.100 90.600 35.200 ;
        RECT 87.000 34.800 90.600 35.100 ;
    END
  END ALU_Out[6]
  PIN ALU_Out[7]
    PORT
      LAYER metal1 ;
        RECT 86.200 58.100 86.600 59.900 ;
        RECT 87.000 58.800 87.400 59.200 ;
        RECT 87.000 58.100 87.300 58.800 ;
        RECT 86.200 57.800 87.300 58.100 ;
        RECT 86.200 55.900 86.600 57.800 ;
        RECT 86.300 54.800 86.600 55.900 ;
        RECT 86.200 51.100 86.600 54.800 ;
      LAYER metal2 ;
        RECT 87.000 58.800 87.400 59.200 ;
        RECT 87.000 58.200 87.300 58.800 ;
        RECT 87.000 57.800 87.400 58.200 ;
      LAYER metal3 ;
        RECT 87.000 58.100 87.400 58.200 ;
        RECT 90.200 58.100 90.600 58.200 ;
        RECT 87.000 57.800 90.600 58.100 ;
    END
  END ALU_Out[7]
  PIN CarryOut
    PORT
      LAYER metal1 ;
        RECT 78.200 66.200 78.600 69.900 ;
        RECT 78.300 65.100 78.600 66.200 ;
        RECT 78.200 61.100 78.600 65.100 ;
      LAYER via1 ;
        RECT 78.200 68.800 78.600 69.200 ;
      LAYER metal2 ;
        RECT 77.400 73.100 77.800 73.200 ;
        RECT 77.400 72.800 78.500 73.100 ;
        RECT 78.200 69.200 78.500 72.800 ;
        RECT 78.200 68.800 78.600 69.200 ;
    END
  END CarryOut
  OBS
      LAYER metal1 ;
        RECT 1.900 68.200 2.300 69.900 ;
        RECT 1.400 67.900 2.300 68.200 ;
        RECT 1.400 61.100 1.800 67.900 ;
        RECT 2.200 67.100 2.600 67.200 ;
        RECT 3.000 67.100 3.400 69.900 ;
        RECT 5.900 68.200 6.300 69.900 ;
        RECT 2.200 66.800 3.400 67.100 ;
        RECT 2.200 65.100 2.600 65.200 ;
        RECT 3.000 65.100 3.400 66.800 ;
        RECT 2.200 64.800 3.400 65.100 ;
        RECT 2.200 64.400 2.600 64.800 ;
        RECT 3.000 61.100 3.400 64.800 ;
        RECT 5.400 67.900 6.300 68.200 ;
        RECT 5.400 67.100 5.800 67.900 ;
        RECT 7.000 67.100 7.400 67.600 ;
        RECT 5.400 66.800 7.400 67.100 ;
        RECT 5.400 61.100 5.800 66.800 ;
        RECT 7.800 61.100 8.200 69.900 ;
        RECT 9.400 66.100 9.800 69.900 ;
        RECT 10.200 68.000 10.600 69.900 ;
        RECT 11.800 68.000 12.200 69.900 ;
        RECT 10.200 67.900 12.200 68.000 ;
        RECT 12.600 67.900 13.000 69.900 ;
        RECT 14.200 68.900 14.600 69.900 ;
        RECT 10.300 67.700 12.100 67.900 ;
        RECT 10.600 67.200 11.000 67.400 ;
        RECT 12.600 67.200 12.900 67.900 ;
        RECT 14.200 67.200 14.500 68.900 ;
        RECT 15.800 68.000 16.200 69.900 ;
        RECT 17.400 68.000 17.800 69.900 ;
        RECT 15.800 67.900 17.800 68.000 ;
        RECT 18.200 67.900 18.600 69.900 ;
        RECT 19.000 67.900 19.400 69.900 ;
        RECT 19.800 68.000 20.200 69.900 ;
        RECT 21.400 68.000 21.800 69.900 ;
        RECT 23.000 68.900 23.400 69.900 ;
        RECT 19.800 67.900 21.800 68.000 ;
        RECT 15.900 67.700 17.700 67.900 ;
        RECT 18.200 67.200 18.500 67.900 ;
        RECT 19.100 67.200 19.400 67.900 ;
        RECT 19.900 67.700 21.700 67.900 ;
        RECT 23.100 67.200 23.400 68.900 ;
        RECT 26.200 67.900 26.600 69.900 ;
        RECT 28.300 68.400 28.700 69.900 ;
        RECT 28.300 67.900 29.000 68.400 ;
        RECT 30.700 68.200 31.100 69.900 ;
        RECT 26.300 67.800 26.600 67.900 ;
        RECT 26.300 67.600 27.200 67.800 ;
        RECT 26.300 67.500 28.400 67.600 ;
        RECT 26.900 67.300 28.400 67.500 ;
        RECT 28.000 67.200 28.400 67.300 ;
        RECT 10.200 66.900 11.000 67.200 ;
        RECT 10.200 66.800 10.600 66.900 ;
        RECT 11.700 66.800 13.000 67.200 ;
        RECT 14.200 66.800 14.600 67.200 ;
        RECT 17.300 66.800 18.600 67.200 ;
        RECT 19.000 66.800 20.300 67.200 ;
        RECT 23.000 66.800 23.400 67.200 ;
        RECT 11.000 66.100 11.400 66.600 ;
        RECT 9.400 65.800 11.400 66.100 ;
        RECT 9.400 61.100 9.800 65.800 ;
        RECT 11.700 65.100 12.000 66.800 ;
        RECT 13.400 65.400 13.800 66.200 ;
        RECT 12.600 65.100 13.000 65.200 ;
        RECT 14.200 65.100 14.500 66.800 ;
        RECT 17.300 65.100 17.600 66.800 ;
        RECT 20.000 66.100 20.300 66.800 ;
        RECT 18.200 65.800 20.300 66.100 ;
        RECT 20.600 65.800 21.000 66.600 ;
        RECT 18.200 65.200 18.500 65.800 ;
        RECT 18.200 65.100 18.600 65.200 ;
        RECT 11.500 64.800 12.000 65.100 ;
        RECT 12.300 64.800 13.000 65.100 ;
        RECT 11.500 64.200 11.900 64.800 ;
        RECT 12.300 64.200 12.600 64.800 ;
        RECT 11.000 63.800 11.900 64.200 ;
        RECT 12.200 63.800 12.600 64.200 ;
        RECT 13.700 64.700 14.600 65.100 ;
        RECT 17.100 64.800 17.600 65.100 ;
        RECT 17.900 64.800 18.600 65.100 ;
        RECT 19.000 65.100 19.400 65.200 ;
        RECT 20.000 65.100 20.300 65.800 ;
        RECT 23.100 65.100 23.400 66.800 ;
        RECT 26.200 66.400 26.600 67.200 ;
        RECT 27.200 66.900 27.600 67.000 ;
        RECT 27.100 66.600 27.600 66.900 ;
        RECT 27.100 66.200 27.400 66.600 ;
        RECT 23.800 65.400 24.200 66.200 ;
        RECT 27.000 65.800 27.400 66.200 ;
        RECT 28.000 65.500 28.300 67.200 ;
        RECT 28.700 66.200 29.000 67.900 ;
        RECT 30.200 68.100 31.100 68.200 ;
        RECT 32.600 68.900 33.000 69.900 ;
        RECT 30.200 67.800 32.100 68.100 ;
        RECT 28.600 65.800 29.000 66.200 ;
        RECT 27.100 65.200 28.300 65.500 ;
        RECT 19.000 64.800 19.700 65.100 ;
        RECT 20.000 64.800 20.500 65.100 ;
        RECT 11.500 61.100 11.900 63.800 ;
        RECT 13.700 62.200 14.100 64.700 ;
        RECT 13.700 61.800 14.600 62.200 ;
        RECT 13.700 61.100 14.100 61.800 ;
        RECT 17.100 61.100 17.500 64.800 ;
        RECT 17.900 64.200 18.200 64.800 ;
        RECT 17.800 63.800 18.200 64.200 ;
        RECT 19.400 64.200 19.700 64.800 ;
        RECT 19.400 63.800 19.800 64.200 ;
        RECT 20.100 61.100 20.500 64.800 ;
        RECT 23.000 64.700 23.900 65.100 ;
        RECT 23.500 62.100 23.900 64.700 ;
        RECT 27.100 63.100 27.400 65.200 ;
        RECT 28.700 65.100 29.000 65.800 ;
        RECT 29.400 65.800 29.800 66.200 ;
        RECT 29.400 65.100 29.700 65.800 ;
        RECT 25.400 62.100 25.800 62.200 ;
        RECT 23.500 61.800 25.800 62.100 ;
        RECT 23.500 61.100 23.900 61.800 ;
        RECT 27.000 61.100 27.400 63.100 ;
        RECT 28.600 64.800 29.700 65.100 ;
        RECT 28.600 61.100 29.000 64.800 ;
        RECT 30.200 61.100 30.600 67.800 ;
        RECT 31.800 67.200 32.100 67.800 ;
        RECT 32.600 67.200 32.900 68.900 ;
        RECT 33.400 67.800 33.800 68.600 ;
        RECT 31.800 66.800 32.200 67.200 ;
        RECT 32.600 66.800 33.000 67.200 ;
        RECT 35.000 67.100 35.400 69.900 ;
        RECT 35.800 68.000 36.200 69.900 ;
        RECT 37.400 68.000 37.800 69.900 ;
        RECT 35.800 67.900 37.800 68.000 ;
        RECT 38.200 67.900 38.600 69.900 ;
        RECT 39.800 68.900 40.200 69.900 ;
        RECT 35.900 67.700 37.700 67.900 ;
        RECT 36.200 67.200 36.600 67.400 ;
        RECT 38.200 67.200 38.500 67.900 ;
        RECT 39.000 67.800 39.400 68.600 ;
        RECT 39.900 67.800 40.200 68.900 ;
        RECT 41.400 67.900 41.800 69.900 ;
        RECT 39.900 67.500 41.100 67.800 ;
        RECT 35.800 67.100 36.600 67.200 ;
        RECT 35.000 66.900 36.600 67.100 ;
        RECT 35.000 66.800 36.200 66.900 ;
        RECT 37.300 66.800 38.600 67.200 ;
        RECT 39.000 67.100 39.400 67.200 ;
        RECT 39.800 67.100 40.300 67.200 ;
        RECT 39.000 66.800 40.300 67.100 ;
        RECT 31.800 65.400 32.200 66.200 ;
        RECT 32.600 65.100 32.900 66.800 ;
        RECT 32.100 64.700 33.000 65.100 ;
        RECT 32.100 61.100 32.500 64.700 ;
        RECT 35.000 61.100 35.400 66.800 ;
        RECT 37.300 65.100 37.600 66.800 ;
        RECT 40.000 66.400 40.400 66.800 ;
        RECT 40.800 66.000 41.100 67.500 ;
        RECT 41.500 66.200 41.800 67.900 ;
        RECT 40.700 65.700 41.100 66.000 ;
        RECT 41.400 65.800 41.800 66.200 ;
        RECT 39.000 65.600 41.100 65.700 ;
        RECT 39.000 65.400 41.000 65.600 ;
        RECT 38.200 65.100 38.600 65.200 ;
        RECT 37.100 64.800 37.600 65.100 ;
        RECT 37.900 64.800 38.600 65.100 ;
        RECT 37.100 61.100 37.500 64.800 ;
        RECT 37.900 64.200 38.200 64.800 ;
        RECT 37.800 63.800 38.200 64.200 ;
        RECT 39.000 61.100 39.400 65.400 ;
        RECT 41.500 65.200 41.800 65.800 ;
        RECT 41.400 65.100 41.800 65.200 ;
        RECT 41.100 64.800 41.800 65.100 ;
        RECT 41.100 61.100 41.500 64.800 ;
        RECT 43.000 61.100 43.400 69.900 ;
        RECT 43.800 67.900 44.200 69.900 ;
        RECT 44.600 68.000 45.000 69.900 ;
        RECT 46.200 68.000 46.600 69.900 ;
        RECT 44.600 67.900 46.600 68.000 ;
        RECT 43.900 67.200 44.200 67.900 ;
        RECT 44.700 67.700 46.500 67.900 ;
        RECT 47.000 67.600 47.400 69.900 ;
        RECT 50.700 67.900 51.500 69.900 ;
        RECT 54.200 68.900 54.600 69.900 ;
        RECT 45.800 67.200 46.200 67.400 ;
        RECT 47.000 67.300 48.100 67.600 ;
        RECT 43.800 66.800 45.100 67.200 ;
        RECT 45.800 66.900 46.600 67.200 ;
        RECT 46.200 66.800 46.600 66.900 ;
        RECT 43.800 66.100 44.200 66.200 ;
        RECT 44.800 66.100 45.100 66.800 ;
        RECT 43.800 65.800 45.100 66.100 ;
        RECT 45.400 65.800 45.800 66.600 ;
        RECT 47.000 65.800 47.400 66.600 ;
        RECT 47.800 65.800 48.100 67.300 ;
        RECT 50.200 66.800 50.600 67.200 ;
        RECT 50.300 66.600 50.600 66.800 ;
        RECT 50.300 66.200 50.700 66.600 ;
        RECT 51.000 66.200 51.300 67.900 ;
        RECT 54.200 67.200 54.500 68.900 ;
        RECT 55.000 67.800 55.400 68.600 ;
        RECT 56.100 68.400 56.500 69.900 ;
        RECT 55.800 67.900 56.500 68.400 ;
        RECT 58.200 67.900 58.600 69.900 ;
        RECT 59.000 68.000 59.400 69.900 ;
        RECT 60.600 68.000 61.000 69.900 ;
        RECT 59.000 67.900 61.000 68.000 ;
        RECT 61.400 67.900 61.800 69.900 ;
        RECT 51.800 67.100 52.200 67.200 ;
        RECT 54.200 67.100 54.600 67.200 ;
        RECT 51.800 66.800 54.600 67.100 ;
        RECT 51.800 66.400 52.200 66.800 ;
        RECT 43.800 65.100 44.200 65.200 ;
        RECT 44.800 65.100 45.100 65.800 ;
        RECT 47.800 65.400 48.400 65.800 ;
        RECT 49.400 65.400 49.800 66.200 ;
        RECT 51.000 65.800 51.400 66.200 ;
        RECT 52.600 66.100 53.000 66.200 ;
        RECT 52.200 65.800 53.000 66.100 ;
        RECT 51.000 65.700 51.300 65.800 ;
        RECT 50.300 65.400 51.300 65.700 ;
        RECT 52.200 65.600 52.600 65.800 ;
        RECT 53.400 65.400 53.800 66.200 ;
        RECT 47.800 65.100 48.100 65.400 ;
        RECT 50.300 65.100 50.600 65.400 ;
        RECT 54.200 65.100 54.500 66.800 ;
        RECT 55.800 66.200 56.100 67.900 ;
        RECT 58.200 67.800 58.500 67.900 ;
        RECT 57.600 67.600 58.500 67.800 ;
        RECT 59.100 67.700 60.900 67.900 ;
        RECT 56.400 67.500 58.500 67.600 ;
        RECT 56.400 67.300 57.900 67.500 ;
        RECT 56.400 67.200 56.800 67.300 ;
        RECT 61.400 67.200 61.700 67.900 ;
        RECT 55.000 66.100 55.400 66.200 ;
        RECT 55.800 66.100 56.200 66.200 ;
        RECT 55.000 65.800 56.200 66.100 ;
        RECT 55.800 65.100 56.100 65.800 ;
        RECT 56.500 65.500 56.800 67.200 ;
        RECT 60.500 66.800 61.800 67.200 ;
        RECT 64.600 67.100 65.000 69.900 ;
        RECT 65.400 68.000 65.800 69.900 ;
        RECT 67.000 68.000 67.400 69.900 ;
        RECT 65.400 67.900 67.400 68.000 ;
        RECT 67.800 67.900 68.200 69.900 ;
        RECT 68.600 67.900 69.000 69.900 ;
        RECT 70.800 68.100 71.600 69.900 ;
        RECT 65.500 67.700 67.300 67.900 ;
        RECT 65.800 67.200 66.200 67.400 ;
        RECT 67.800 67.200 68.100 67.900 ;
        RECT 68.600 67.600 69.700 67.900 ;
        RECT 69.300 67.500 69.700 67.600 ;
        RECT 65.400 67.100 66.200 67.200 ;
        RECT 64.600 66.900 66.200 67.100 ;
        RECT 64.600 66.800 65.800 66.900 ;
        RECT 66.900 66.800 68.200 67.200 ;
        RECT 56.500 65.200 57.700 65.500 ;
        RECT 43.800 64.800 44.500 65.100 ;
        RECT 44.800 64.800 45.300 65.100 ;
        RECT 44.200 64.200 44.500 64.800 ;
        RECT 44.200 63.800 44.600 64.200 ;
        RECT 44.900 61.100 45.300 64.800 ;
        RECT 47.000 64.800 48.100 65.100 ;
        RECT 47.000 61.100 47.400 64.800 ;
        RECT 49.400 61.400 49.800 65.100 ;
        RECT 50.200 61.700 50.600 65.100 ;
        RECT 51.000 64.800 53.000 65.100 ;
        RECT 51.000 61.400 51.400 64.800 ;
        RECT 49.400 61.100 51.400 61.400 ;
        RECT 52.600 61.100 53.000 64.800 ;
        RECT 53.700 64.700 54.600 65.100 ;
        RECT 53.700 61.100 54.100 64.700 ;
        RECT 55.800 61.100 56.200 65.100 ;
        RECT 57.400 63.100 57.700 65.200 ;
        RECT 60.500 65.100 60.800 66.800 ;
        RECT 61.400 65.100 61.800 65.200 ;
        RECT 60.300 64.800 60.800 65.100 ;
        RECT 61.100 64.800 61.800 65.100 ;
        RECT 57.400 61.100 57.800 63.100 ;
        RECT 60.300 62.200 60.700 64.800 ;
        RECT 61.100 64.200 61.400 64.800 ;
        RECT 61.000 63.800 61.800 64.200 ;
        RECT 59.800 61.800 60.700 62.200 ;
        RECT 60.300 61.100 60.700 61.800 ;
        RECT 64.600 61.100 65.000 66.800 ;
        RECT 66.900 65.100 67.200 66.800 ;
        RECT 70.600 66.700 71.000 67.100 ;
        RECT 70.600 66.400 70.900 66.700 ;
        RECT 69.600 66.100 70.900 66.400 ;
        RECT 71.300 66.400 71.600 68.100 ;
        RECT 73.400 67.900 73.800 69.900 ;
        RECT 74.500 68.200 74.900 69.900 ;
        RECT 74.500 67.900 75.400 68.200 ;
        RECT 72.600 67.600 73.800 67.900 ;
        RECT 72.600 67.500 73.000 67.600 ;
        RECT 71.300 66.200 71.800 66.400 ;
        RECT 71.300 66.100 72.200 66.200 ;
        RECT 69.600 66.000 70.000 66.100 ;
        RECT 71.500 65.800 72.200 66.100 ;
        RECT 70.700 65.700 71.100 65.800 ;
        RECT 69.400 65.400 71.100 65.700 ;
        RECT 67.800 65.100 68.200 65.200 ;
        RECT 69.400 65.100 69.700 65.400 ;
        RECT 71.500 65.100 71.800 65.800 ;
        RECT 66.700 64.800 67.200 65.100 ;
        RECT 67.500 64.800 68.200 65.100 ;
        RECT 68.600 64.800 69.700 65.100 ;
        RECT 66.700 61.100 67.100 64.800 ;
        RECT 67.500 64.200 67.800 64.800 ;
        RECT 67.400 63.800 67.800 64.200 ;
        RECT 68.600 61.100 69.000 64.800 ;
        RECT 69.300 64.700 69.700 64.800 ;
        RECT 70.800 64.800 71.800 65.100 ;
        RECT 72.600 64.800 73.800 65.100 ;
        RECT 70.800 61.100 71.600 64.800 ;
        RECT 72.600 64.700 73.000 64.800 ;
        RECT 73.400 61.100 73.800 64.800 ;
        RECT 74.200 64.400 74.600 65.200 ;
        RECT 75.000 61.100 75.400 67.900 ;
        RECT 76.600 67.600 77.000 69.900 ;
        RECT 79.800 68.900 80.200 69.900 ;
        RECT 75.800 66.800 76.200 67.600 ;
        RECT 76.600 67.300 77.700 67.600 ;
        RECT 76.600 65.800 77.000 66.600 ;
        RECT 77.400 65.800 77.700 67.300 ;
        RECT 79.900 67.200 80.200 68.900 ;
        RECT 82.700 68.200 83.100 69.900 ;
        RECT 82.200 67.900 83.100 68.200 ;
        RECT 79.800 66.800 80.200 67.200 ;
        RECT 81.400 67.100 81.800 67.600 ;
        RECT 77.400 65.400 78.000 65.800 ;
        RECT 77.400 65.100 77.700 65.400 ;
        RECT 79.900 65.100 80.200 66.800 ;
        RECT 80.600 66.800 81.800 67.100 ;
        RECT 80.600 66.200 80.900 66.800 ;
        RECT 80.600 65.400 81.000 66.200 ;
        RECT 76.600 64.800 77.700 65.100 ;
        RECT 76.600 61.100 77.000 64.800 ;
        RECT 79.800 64.700 80.700 65.100 ;
        RECT 80.300 62.200 80.700 64.700 ;
        RECT 80.300 61.800 81.000 62.200 ;
        RECT 80.300 61.100 80.700 61.800 ;
        RECT 82.200 61.100 82.600 67.900 ;
        RECT 83.000 65.100 83.400 65.200 ;
        RECT 83.800 65.100 84.200 69.900 ;
        RECT 83.000 64.800 84.200 65.100 ;
        RECT 83.000 64.400 83.400 64.800 ;
        RECT 83.800 61.100 84.200 64.800 ;
        RECT 1.400 55.100 1.800 59.900 ;
        RECT 3.500 56.300 3.900 59.900 ;
        RECT 3.000 55.900 3.900 56.300 ;
        RECT 2.200 55.100 2.600 55.200 ;
        RECT 1.400 54.800 2.600 55.100 ;
        RECT 1.400 51.100 1.800 54.800 ;
        RECT 3.100 54.200 3.400 55.900 ;
        RECT 4.600 55.800 5.000 56.600 ;
        RECT 3.800 55.100 4.200 55.600 ;
        RECT 4.600 55.100 4.900 55.800 ;
        RECT 3.800 54.800 4.900 55.100 ;
        RECT 3.000 53.800 3.400 54.200 ;
        RECT 3.100 52.200 3.400 53.800 ;
        RECT 5.400 53.100 5.800 59.900 ;
        RECT 7.000 55.900 7.400 59.900 ;
        RECT 7.800 56.200 8.200 59.900 ;
        RECT 9.400 56.200 9.800 59.900 ;
        RECT 7.800 55.900 9.800 56.200 ;
        RECT 10.500 56.300 10.900 59.900 ;
        RECT 10.500 55.900 11.400 56.300 ;
        RECT 13.400 56.100 13.800 59.900 ;
        RECT 14.200 56.100 14.600 56.600 ;
        RECT 7.100 55.200 7.400 55.900 ;
        RECT 9.000 55.200 9.400 55.400 ;
        RECT 7.000 54.900 8.200 55.200 ;
        RECT 9.000 54.900 9.800 55.200 ;
        RECT 7.000 54.800 7.400 54.900 ;
        RECT 3.000 51.100 3.400 52.200 ;
        RECT 4.900 52.800 5.800 53.100 ;
        RECT 7.000 52.800 7.400 53.200 ;
        RECT 7.900 53.100 8.200 54.900 ;
        RECT 9.400 54.800 9.800 54.900 ;
        RECT 10.200 54.800 10.600 55.600 ;
        RECT 8.600 53.800 9.000 54.600 ;
        RECT 11.000 54.200 11.300 55.900 ;
        RECT 13.400 55.800 14.600 56.100 ;
        RECT 15.000 56.100 15.400 59.900 ;
        RECT 17.000 56.800 17.400 57.200 ;
        RECT 17.000 56.200 17.300 56.800 ;
        RECT 17.700 56.200 18.100 59.900 ;
        RECT 16.600 56.100 17.300 56.200 ;
        RECT 15.000 55.900 17.300 56.100 ;
        RECT 17.600 55.900 18.100 56.200 ;
        RECT 19.800 55.900 20.200 59.900 ;
        RECT 20.600 56.200 21.000 59.900 ;
        RECT 22.200 56.200 22.600 59.900 ;
        RECT 20.600 55.900 22.600 56.200 ;
        RECT 25.900 56.200 26.300 59.900 ;
        RECT 26.600 56.800 27.000 57.200 ;
        RECT 26.700 56.200 27.000 56.800 ;
        RECT 27.800 56.200 28.200 59.900 ;
        RECT 28.700 56.200 29.100 56.300 ;
        RECT 25.900 55.900 26.400 56.200 ;
        RECT 26.700 55.900 27.400 56.200 ;
        RECT 27.800 55.900 29.100 56.200 ;
        RECT 30.000 55.900 30.800 59.900 ;
        RECT 31.800 56.200 32.200 56.300 ;
        RECT 32.600 56.200 33.000 59.900 ;
        RECT 31.800 55.900 33.000 56.200 ;
        RECT 33.400 59.600 35.400 59.900 ;
        RECT 33.400 55.900 33.800 59.600 ;
        RECT 34.200 55.900 34.600 59.300 ;
        RECT 35.000 56.200 35.400 59.600 ;
        RECT 36.600 56.200 37.000 59.900 ;
        RECT 35.000 55.900 37.000 56.200 ;
        RECT 15.000 55.800 17.000 55.900 ;
        RECT 11.000 53.800 11.400 54.200 ;
        RECT 13.400 54.100 13.800 55.800 ;
        RECT 11.800 53.800 13.800 54.100 ;
        RECT 14.200 54.800 14.600 55.200 ;
        RECT 14.200 54.100 14.500 54.800 ;
        RECT 15.000 54.100 15.400 55.800 ;
        RECT 17.600 54.200 17.900 55.900 ;
        RECT 19.900 55.200 20.200 55.900 ;
        RECT 21.800 55.200 22.200 55.400 ;
        RECT 18.200 54.400 18.600 55.200 ;
        RECT 19.800 54.900 21.000 55.200 ;
        RECT 21.800 54.900 22.600 55.200 ;
        RECT 19.800 54.800 20.200 54.900 ;
        RECT 14.200 53.800 15.400 54.100 ;
        RECT 16.600 53.800 17.900 54.200 ;
        RECT 19.000 54.100 19.400 54.200 ;
        RECT 18.600 53.800 19.400 54.100 ;
        RECT 4.900 52.200 5.300 52.800 ;
        RECT 7.100 52.400 7.500 52.800 ;
        RECT 4.900 51.800 5.800 52.200 ;
        RECT 4.900 51.100 5.300 51.800 ;
        RECT 7.800 51.100 8.200 53.100 ;
        RECT 11.000 52.200 11.300 53.800 ;
        RECT 11.800 53.200 12.100 53.800 ;
        RECT 11.800 52.400 12.200 53.200 ;
        RECT 11.000 51.100 11.400 52.200 ;
        RECT 13.400 51.100 13.800 53.800 ;
        RECT 15.000 53.100 15.400 53.800 ;
        RECT 16.700 53.100 17.000 53.800 ;
        RECT 18.600 53.600 19.000 53.800 ;
        RECT 17.500 53.100 19.300 53.300 ;
        RECT 14.500 52.800 15.400 53.100 ;
        RECT 14.500 51.100 14.900 52.800 ;
        RECT 16.600 51.100 17.000 53.100 ;
        RECT 17.400 53.000 19.400 53.100 ;
        RECT 17.400 51.100 17.800 53.000 ;
        RECT 19.000 51.100 19.400 53.000 ;
        RECT 19.800 52.800 20.200 53.200 ;
        RECT 20.700 53.100 21.000 54.900 ;
        RECT 22.200 54.800 22.600 54.900 ;
        RECT 21.400 54.100 21.800 54.600 ;
        RECT 26.100 54.200 26.400 55.900 ;
        RECT 27.000 55.800 27.400 55.900 ;
        RECT 29.300 55.200 29.700 55.300 ;
        RECT 30.300 55.200 30.600 55.900 ;
        RECT 34.300 55.600 34.600 55.900 ;
        RECT 34.300 55.300 35.300 55.600 ;
        RECT 28.900 54.900 29.700 55.200 ;
        RECT 28.900 54.800 29.300 54.900 ;
        RECT 30.200 54.800 30.600 55.200 ;
        RECT 35.000 55.200 35.300 55.300 ;
        RECT 36.200 55.200 36.600 55.400 ;
        RECT 35.000 54.800 35.400 55.200 ;
        RECT 36.200 54.900 37.000 55.200 ;
        RECT 36.600 54.800 37.000 54.900 ;
        RECT 38.200 55.100 38.600 59.900 ;
        RECT 39.000 56.100 39.400 56.600 ;
        RECT 39.800 56.100 40.200 59.900 ;
        RECT 39.000 55.800 40.200 56.100 ;
        RECT 38.200 54.800 39.300 55.100 ;
        RECT 30.300 54.200 30.600 54.800 ;
        RECT 34.300 54.400 34.700 54.800 ;
        RECT 34.300 54.200 34.600 54.400 ;
        RECT 23.000 54.100 23.400 54.200 ;
        RECT 21.400 53.800 23.400 54.100 ;
        RECT 26.100 53.800 27.400 54.200 ;
        RECT 30.300 53.900 30.800 54.200 ;
        RECT 24.700 53.100 26.500 53.300 ;
        RECT 27.000 53.100 27.300 53.800 ;
        RECT 28.700 53.400 29.100 53.500 ;
        RECT 27.800 53.100 29.100 53.400 ;
        RECT 29.400 53.200 30.200 53.600 ;
        RECT 19.900 52.400 20.300 52.800 ;
        RECT 20.600 51.100 21.000 53.100 ;
        RECT 24.600 53.000 26.600 53.100 ;
        RECT 24.600 51.100 25.000 53.000 ;
        RECT 26.200 51.100 26.600 53.000 ;
        RECT 27.000 51.100 27.400 53.100 ;
        RECT 27.800 51.100 28.200 53.100 ;
        RECT 30.500 52.900 30.800 53.900 ;
        RECT 31.200 53.800 31.600 54.200 ;
        RECT 34.200 53.800 34.600 54.200 ;
        RECT 31.200 53.600 31.500 53.800 ;
        RECT 31.100 53.200 31.500 53.600 ;
        RECT 31.800 53.400 32.200 53.500 ;
        RECT 31.800 53.100 33.000 53.400 ;
        RECT 35.000 53.100 35.300 54.800 ;
        RECT 35.800 53.800 36.200 54.600 ;
        RECT 38.200 53.100 38.600 54.800 ;
        RECT 39.000 54.200 39.300 54.800 ;
        RECT 39.000 53.800 39.400 54.200 ;
        RECT 39.800 54.100 40.200 55.800 ;
        RECT 41.400 54.100 41.800 54.200 ;
        RECT 39.800 53.800 41.800 54.100 ;
        RECT 30.000 52.200 30.800 52.900 ;
        RECT 29.400 51.800 30.800 52.200 ;
        RECT 30.000 51.100 30.800 51.800 ;
        RECT 32.600 51.100 33.000 53.100 ;
        RECT 34.700 51.100 35.500 53.100 ;
        RECT 38.200 52.800 39.100 53.100 ;
        RECT 38.700 51.100 39.100 52.800 ;
        RECT 39.800 51.100 40.200 53.800 ;
        RECT 41.400 53.400 41.800 53.800 ;
        RECT 42.200 53.100 42.600 59.900 ;
        RECT 43.000 56.100 43.400 56.600 ;
        RECT 43.800 56.100 44.200 56.200 ;
        RECT 43.000 55.800 44.200 56.100 ;
        RECT 44.600 53.100 45.000 59.900 ;
        RECT 45.400 55.800 45.800 56.600 ;
        RECT 47.500 56.300 47.900 59.900 ;
        RECT 47.000 55.900 47.900 56.300 ;
        RECT 48.900 56.300 49.300 59.900 ;
        RECT 48.900 55.900 49.800 56.300 ;
        RECT 51.800 56.100 52.200 59.900 ;
        RECT 52.600 56.800 53.000 57.200 ;
        RECT 52.600 56.100 52.900 56.800 ;
        RECT 47.100 54.200 47.400 55.900 ;
        RECT 47.800 55.100 48.200 55.600 ;
        RECT 48.600 55.100 49.000 55.600 ;
        RECT 47.800 54.800 49.000 55.100 ;
        RECT 47.000 53.800 47.400 54.200 ;
        RECT 42.200 52.800 43.100 53.100 ;
        RECT 44.600 52.800 45.500 53.100 ;
        RECT 42.700 52.200 43.100 52.800 ;
        RECT 42.200 51.800 43.100 52.200 ;
        RECT 42.700 51.100 43.100 51.800 ;
        RECT 45.100 52.200 45.500 52.800 ;
        RECT 47.100 52.200 47.400 53.800 ;
        RECT 45.100 51.800 45.800 52.200 ;
        RECT 45.100 51.100 45.500 51.800 ;
        RECT 47.000 51.100 47.400 52.200 ;
        RECT 49.400 54.200 49.700 55.900 ;
        RECT 51.800 55.800 52.900 56.100 ;
        RECT 49.400 53.800 49.800 54.200 ;
        RECT 49.400 52.200 49.700 53.800 ;
        RECT 50.200 52.400 50.600 53.200 ;
        RECT 49.400 51.100 49.800 52.200 ;
        RECT 51.800 51.100 52.200 55.800 ;
        RECT 52.600 55.100 53.000 55.200 ;
        RECT 53.400 55.100 53.800 59.900 ;
        RECT 52.600 54.800 53.800 55.100 ;
        RECT 54.200 55.800 54.600 56.600 ;
        RECT 55.300 56.300 55.700 59.900 ;
        RECT 55.300 55.900 56.200 56.300 ;
        RECT 54.200 55.100 54.500 55.800 ;
        RECT 55.000 55.100 55.400 55.600 ;
        RECT 54.200 54.800 55.400 55.100 ;
        RECT 55.800 55.100 56.100 55.900 ;
        RECT 55.800 54.800 57.700 55.100 ;
        RECT 53.400 53.100 53.800 54.800 ;
        RECT 55.800 54.200 56.100 54.800 ;
        RECT 57.400 54.200 57.700 54.800 ;
        RECT 55.800 53.800 56.200 54.200 ;
        RECT 53.400 52.800 54.300 53.100 ;
        RECT 53.900 51.100 54.300 52.800 ;
        RECT 55.800 52.100 56.100 53.800 ;
        RECT 57.400 53.400 57.800 54.200 ;
        RECT 55.800 51.100 56.200 52.100 ;
        RECT 58.200 51.100 58.600 59.900 ;
        RECT 59.000 53.400 59.400 54.200 ;
        RECT 59.800 53.100 60.200 59.900 ;
        RECT 63.800 57.900 64.200 59.900 ;
        RECT 63.900 57.800 64.200 57.900 ;
        RECT 65.400 57.900 65.800 59.900 ;
        RECT 65.400 57.800 65.700 57.900 ;
        RECT 63.900 57.500 65.700 57.800 ;
        RECT 60.600 55.800 61.000 56.600 ;
        RECT 64.600 56.400 65.000 57.200 ;
        RECT 65.400 56.200 65.700 57.500 ;
        RECT 66.200 56.200 66.600 59.900 ;
        RECT 67.800 59.600 69.800 59.900 ;
        RECT 67.800 56.200 68.200 59.600 ;
        RECT 63.000 55.400 63.400 56.200 ;
        RECT 65.400 55.800 65.800 56.200 ;
        RECT 66.200 55.900 68.200 56.200 ;
        RECT 68.600 55.900 69.000 59.300 ;
        RECT 69.400 55.900 69.800 59.600 ;
        RECT 63.800 54.800 64.600 55.200 ;
        RECT 65.400 54.200 65.700 55.800 ;
        RECT 68.600 55.600 68.900 55.900 ;
        RECT 66.600 55.200 67.000 55.400 ;
        RECT 67.900 55.300 68.900 55.600 ;
        RECT 67.900 55.200 68.200 55.300 ;
        RECT 64.900 54.100 65.700 54.200 ;
        RECT 64.800 53.900 65.700 54.100 ;
        RECT 66.200 54.900 67.000 55.200 ;
        RECT 66.200 54.800 66.600 54.900 ;
        RECT 67.800 54.800 68.200 55.200 ;
        RECT 69.400 55.100 69.800 55.600 ;
        RECT 70.200 55.100 70.600 59.900 ;
        RECT 72.900 59.200 73.300 59.900 ;
        RECT 72.900 58.800 73.800 59.200 ;
        RECT 72.200 56.800 72.600 57.200 ;
        RECT 72.200 56.200 72.500 56.800 ;
        RECT 72.900 56.200 73.300 58.800 ;
        RECT 71.800 55.900 72.500 56.200 ;
        RECT 72.800 55.900 73.300 56.200 ;
        RECT 75.000 56.200 75.400 59.900 ;
        RECT 76.600 56.200 77.000 59.900 ;
        RECT 75.000 55.900 77.000 56.200 ;
        RECT 77.400 55.900 77.800 59.900 ;
        RECT 78.200 55.900 78.600 59.900 ;
        RECT 79.000 56.200 79.400 59.900 ;
        RECT 80.600 56.200 81.000 59.900 ;
        RECT 82.200 57.900 82.600 59.900 ;
        RECT 82.300 57.800 82.600 57.900 ;
        RECT 83.800 57.900 84.200 59.900 ;
        RECT 83.800 57.800 84.100 57.900 ;
        RECT 82.300 57.500 84.100 57.800 ;
        RECT 79.000 55.900 81.000 56.200 ;
        RECT 71.800 55.800 72.200 55.900 ;
        RECT 69.400 54.800 70.600 55.100 ;
        RECT 66.200 54.200 66.500 54.800 ;
        RECT 64.800 53.200 65.200 53.900 ;
        RECT 66.200 53.800 66.600 54.200 ;
        RECT 67.000 53.800 67.400 54.600 ;
        RECT 59.800 52.800 60.700 53.100 ;
        RECT 60.300 52.100 60.700 52.800 ;
        RECT 62.200 52.800 62.600 53.200 ;
        RECT 64.800 52.800 65.800 53.200 ;
        RECT 67.900 53.100 68.200 54.800 ;
        RECT 68.500 54.400 68.900 54.800 ;
        RECT 68.600 54.200 68.900 54.400 ;
        RECT 68.600 54.100 69.000 54.200 ;
        RECT 69.400 54.100 69.800 54.200 ;
        RECT 68.600 53.800 69.800 54.100 ;
        RECT 62.200 52.100 62.500 52.800 ;
        RECT 60.300 51.800 62.500 52.100 ;
        RECT 60.300 51.100 60.700 51.800 ;
        RECT 64.800 51.100 65.200 52.800 ;
        RECT 67.700 51.100 68.500 53.100 ;
        RECT 70.200 51.100 70.600 54.800 ;
        RECT 72.800 54.200 73.100 55.900 ;
        RECT 75.400 55.200 75.800 55.400 ;
        RECT 77.400 55.200 77.700 55.900 ;
        RECT 78.300 55.200 78.600 55.900 ;
        RECT 80.200 55.200 80.600 55.400 ;
        RECT 73.400 54.400 73.800 55.200 ;
        RECT 75.000 54.900 75.800 55.200 ;
        RECT 76.600 54.900 77.800 55.200 ;
        RECT 75.000 54.800 75.400 54.900 ;
        RECT 71.000 53.400 71.400 54.200 ;
        RECT 71.800 53.800 73.100 54.200 ;
        RECT 74.200 54.100 74.600 54.200 ;
        RECT 73.800 53.800 74.600 54.100 ;
        RECT 75.800 53.800 76.200 54.600 ;
        RECT 76.600 54.100 76.900 54.900 ;
        RECT 77.400 54.800 77.800 54.900 ;
        RECT 78.200 54.900 79.400 55.200 ;
        RECT 80.200 54.900 81.000 55.200 ;
        RECT 78.200 54.800 78.600 54.900 ;
        RECT 77.400 54.100 77.800 54.200 ;
        RECT 76.600 53.800 77.800 54.100 ;
        RECT 71.900 53.100 72.200 53.800 ;
        RECT 73.800 53.600 74.200 53.800 ;
        RECT 72.700 53.100 74.500 53.300 ;
        RECT 76.600 53.100 76.900 53.800 ;
        RECT 71.800 51.100 72.200 53.100 ;
        RECT 72.600 53.000 74.600 53.100 ;
        RECT 72.600 51.100 73.000 53.000 ;
        RECT 74.200 51.100 74.600 53.000 ;
        RECT 76.600 51.100 77.000 53.100 ;
        RECT 77.400 52.800 77.800 53.200 ;
        RECT 78.200 52.800 78.600 53.200 ;
        RECT 79.100 53.100 79.400 54.900 ;
        RECT 80.600 54.800 81.000 54.900 ;
        RECT 81.400 54.800 81.800 56.200 ;
        RECT 83.000 55.800 83.400 57.200 ;
        RECT 83.800 56.200 84.100 57.500 ;
        RECT 84.600 56.200 85.000 59.900 ;
        RECT 83.800 55.800 84.200 56.200 ;
        RECT 84.600 55.900 85.700 56.200 ;
        RECT 82.200 54.800 83.000 55.200 ;
        RECT 79.800 53.800 80.200 54.600 ;
        RECT 83.800 54.200 84.100 55.800 ;
        RECT 85.400 55.600 85.700 55.900 ;
        RECT 85.400 55.200 86.000 55.600 ;
        RECT 84.600 54.400 85.000 55.200 ;
        RECT 83.300 54.100 84.100 54.200 ;
        RECT 82.200 53.900 84.100 54.100 ;
        RECT 82.200 53.800 83.600 53.900 ;
        RECT 77.300 52.400 77.700 52.800 ;
        RECT 78.300 52.400 78.700 52.800 ;
        RECT 79.000 51.100 79.400 53.100 ;
        RECT 82.200 53.200 82.500 53.800 ;
        RECT 82.200 52.800 82.600 53.200 ;
        RECT 83.200 51.100 83.600 53.800 ;
        RECT 85.400 53.700 85.700 55.200 ;
        RECT 84.600 53.400 85.700 53.700 ;
        RECT 84.600 51.100 85.000 53.400 ;
        RECT 2.200 47.600 2.600 49.900 ;
        RECT 3.100 48.200 3.500 48.600 ;
        RECT 3.000 47.800 3.400 48.200 ;
        RECT 3.800 47.900 4.200 49.900 ;
        RECT 6.200 47.900 6.600 49.900 ;
        RECT 7.000 48.000 7.400 49.900 ;
        RECT 8.600 48.000 9.000 49.900 ;
        RECT 7.000 47.900 9.000 48.000 ;
        RECT 9.400 47.900 9.800 49.900 ;
        RECT 10.200 48.000 10.600 49.900 ;
        RECT 11.800 48.000 12.200 49.900 ;
        RECT 12.900 49.200 13.300 49.900 ;
        RECT 12.600 48.800 13.300 49.200 ;
        RECT 12.900 48.400 13.300 48.800 ;
        RECT 10.200 47.900 12.200 48.000 ;
        RECT 12.600 47.900 13.300 48.400 ;
        RECT 15.000 47.900 15.400 49.900 ;
        RECT 15.800 48.000 16.200 49.900 ;
        RECT 17.400 48.000 17.800 49.900 ;
        RECT 15.800 47.900 17.800 48.000 ;
        RECT 18.200 47.900 18.600 49.900 ;
        RECT 19.100 48.200 19.500 48.600 ;
        RECT 1.500 47.300 2.600 47.600 ;
        RECT 1.500 45.800 1.800 47.300 ;
        RECT 2.200 45.800 2.600 46.600 ;
        RECT 3.900 46.200 4.200 47.900 ;
        RECT 6.300 47.200 6.600 47.900 ;
        RECT 7.100 47.700 8.900 47.900 ;
        RECT 8.200 47.200 8.600 47.400 ;
        RECT 9.500 47.200 9.800 47.900 ;
        RECT 10.300 47.700 12.100 47.900 ;
        RECT 11.400 47.200 11.800 47.400 ;
        RECT 4.600 46.400 5.000 47.200 ;
        RECT 6.200 46.800 7.500 47.200 ;
        RECT 8.200 46.900 9.000 47.200 ;
        RECT 8.600 46.800 9.000 46.900 ;
        RECT 9.400 46.800 10.700 47.200 ;
        RECT 11.400 46.900 12.200 47.200 ;
        RECT 11.800 46.800 12.200 46.900 ;
        RECT 3.000 46.100 3.400 46.200 ;
        RECT 3.800 46.100 4.200 46.200 ;
        RECT 5.400 46.100 5.800 46.200 ;
        RECT 3.000 45.800 4.200 46.100 ;
        RECT 5.000 45.800 5.800 46.100 ;
        RECT 6.200 46.100 6.600 46.200 ;
        RECT 7.200 46.100 7.500 46.800 ;
        RECT 6.200 45.800 7.500 46.100 ;
        RECT 7.800 46.100 8.200 46.600 ;
        RECT 10.400 46.100 10.700 46.800 ;
        RECT 7.800 45.800 10.700 46.100 ;
        RECT 11.000 45.800 11.400 46.600 ;
        RECT 12.600 46.200 12.900 47.900 ;
        RECT 15.000 47.800 15.300 47.900 ;
        RECT 14.400 47.600 15.300 47.800 ;
        RECT 15.900 47.700 17.700 47.900 ;
        RECT 13.200 47.500 15.300 47.600 ;
        RECT 13.200 47.300 14.700 47.500 ;
        RECT 13.200 47.200 13.600 47.300 ;
        RECT 16.200 47.200 16.600 47.400 ;
        RECT 18.200 47.200 18.500 47.900 ;
        RECT 19.000 47.800 19.400 48.200 ;
        RECT 19.800 47.900 20.200 49.900 ;
        RECT 12.600 45.800 13.000 46.200 ;
        RECT 1.200 45.400 1.800 45.800 ;
        RECT 1.500 45.100 1.800 45.400 ;
        RECT 3.100 45.100 3.400 45.800 ;
        RECT 5.000 45.600 5.400 45.800 ;
        RECT 6.200 45.100 6.600 45.200 ;
        RECT 7.200 45.100 7.500 45.800 ;
        RECT 9.400 45.100 9.800 45.200 ;
        RECT 10.400 45.100 10.700 45.800 ;
        RECT 12.600 45.100 12.900 45.800 ;
        RECT 13.300 45.500 13.600 47.200 ;
        RECT 14.000 46.900 14.400 47.000 ;
        RECT 14.000 46.600 14.500 46.900 ;
        RECT 14.200 46.200 14.500 46.600 ;
        RECT 15.000 46.400 15.400 47.200 ;
        RECT 15.800 46.900 16.600 47.200 ;
        RECT 15.800 46.800 16.200 46.900 ;
        RECT 17.300 46.800 18.600 47.200 ;
        RECT 14.200 45.800 14.600 46.200 ;
        RECT 16.600 45.800 17.000 46.600 ;
        RECT 13.300 45.200 14.500 45.500 ;
        RECT 1.500 44.800 2.600 45.100 ;
        RECT 2.200 41.100 2.600 44.800 ;
        RECT 3.000 41.100 3.400 45.100 ;
        RECT 3.800 44.800 5.800 45.100 ;
        RECT 6.200 44.800 6.900 45.100 ;
        RECT 7.200 44.800 7.700 45.100 ;
        RECT 9.400 44.800 10.100 45.100 ;
        RECT 10.400 44.800 10.900 45.100 ;
        RECT 3.800 41.100 4.200 44.800 ;
        RECT 5.400 41.100 5.800 44.800 ;
        RECT 6.600 44.200 6.900 44.800 ;
        RECT 6.600 43.800 7.000 44.200 ;
        RECT 7.300 41.100 7.700 44.800 ;
        RECT 9.800 44.200 10.100 44.800 ;
        RECT 9.800 43.800 10.200 44.200 ;
        RECT 10.500 41.100 10.900 44.800 ;
        RECT 12.600 41.100 13.000 45.100 ;
        RECT 14.200 43.100 14.500 45.200 ;
        RECT 17.300 45.100 17.600 46.800 ;
        RECT 19.000 46.100 19.400 46.200 ;
        RECT 19.900 46.100 20.200 47.900 ;
        RECT 20.600 46.400 21.000 47.200 ;
        RECT 21.400 47.100 21.800 47.200 ;
        RECT 22.200 47.100 22.600 49.900 ;
        RECT 25.400 48.000 25.800 49.900 ;
        RECT 27.000 48.000 27.400 49.900 ;
        RECT 25.400 47.900 27.400 48.000 ;
        RECT 27.800 48.100 28.200 49.900 ;
        RECT 29.400 48.900 29.800 49.900 ;
        RECT 28.600 48.100 29.000 48.600 ;
        RECT 25.500 47.700 27.300 47.900 ;
        RECT 27.800 47.800 29.000 48.100 ;
        RECT 21.400 46.800 22.600 47.100 ;
        RECT 23.000 46.800 23.400 47.600 ;
        RECT 25.800 47.200 26.200 47.400 ;
        RECT 27.800 47.200 28.100 47.800 ;
        RECT 29.500 47.200 29.800 48.900 ;
        RECT 31.000 48.000 31.400 49.900 ;
        RECT 32.600 48.000 33.000 49.900 ;
        RECT 31.000 47.900 33.000 48.000 ;
        RECT 33.400 47.900 33.800 49.900 ;
        RECT 35.500 47.900 36.300 49.900 ;
        RECT 31.100 47.700 32.900 47.900 ;
        RECT 31.400 47.200 31.800 47.400 ;
        RECT 33.400 47.200 33.700 47.900 ;
        RECT 25.400 46.900 26.200 47.200 ;
        RECT 25.400 46.800 25.800 46.900 ;
        RECT 26.900 46.800 28.200 47.200 ;
        RECT 29.400 47.100 29.800 47.200 ;
        RECT 28.600 46.800 29.800 47.100 ;
        RECT 31.000 46.900 31.800 47.200 ;
        RECT 31.000 46.800 31.400 46.900 ;
        RECT 32.500 46.800 33.800 47.200 ;
        RECT 35.000 46.800 35.400 47.200 ;
        RECT 21.400 46.100 21.800 46.200 ;
        RECT 22.200 46.100 22.600 46.800 ;
        RECT 26.200 46.100 26.600 46.600 ;
        RECT 19.000 45.800 20.200 46.100 ;
        RECT 21.000 45.800 26.600 46.100 ;
        RECT 18.200 45.100 18.600 45.200 ;
        RECT 19.100 45.100 19.400 45.800 ;
        RECT 21.000 45.600 21.400 45.800 ;
        RECT 17.100 44.800 17.600 45.100 ;
        RECT 17.900 44.800 19.400 45.100 ;
        RECT 14.200 41.100 14.600 43.100 ;
        RECT 17.100 41.100 17.500 44.800 ;
        RECT 17.900 44.200 18.200 44.800 ;
        RECT 17.800 43.800 18.200 44.200 ;
        RECT 19.000 41.100 19.400 44.800 ;
        RECT 19.800 44.800 21.800 45.100 ;
        RECT 19.800 41.100 20.200 44.800 ;
        RECT 21.400 41.100 21.800 44.800 ;
        RECT 22.200 41.100 22.600 45.800 ;
        RECT 26.900 45.100 27.200 46.800 ;
        RECT 28.600 46.200 28.900 46.800 ;
        RECT 28.600 45.800 29.000 46.200 ;
        RECT 27.800 45.100 28.200 45.200 ;
        RECT 29.500 45.100 29.800 46.800 ;
        RECT 30.200 45.400 30.600 46.200 ;
        RECT 31.000 46.100 31.400 46.200 ;
        RECT 31.800 46.100 32.200 46.600 ;
        RECT 31.000 45.800 32.200 46.100 ;
        RECT 32.500 45.200 32.800 46.800 ;
        RECT 35.100 46.600 35.400 46.800 ;
        RECT 35.100 46.200 35.500 46.600 ;
        RECT 35.800 46.200 36.100 47.900 ;
        RECT 36.600 46.400 37.000 47.200 ;
        RECT 35.800 45.800 36.200 46.200 ;
        RECT 37.400 46.100 37.800 46.200 ;
        RECT 37.000 45.800 37.800 46.100 ;
        RECT 35.800 45.700 36.100 45.800 ;
        RECT 35.100 45.400 36.100 45.700 ;
        RECT 37.000 45.600 37.400 45.800 ;
        RECT 35.100 45.200 35.400 45.400 ;
        RECT 26.700 44.800 27.200 45.100 ;
        RECT 27.500 44.800 28.200 45.100 ;
        RECT 26.700 41.100 27.100 44.800 ;
        RECT 27.500 44.200 27.800 44.800 ;
        RECT 29.400 44.700 30.300 45.100 ;
        RECT 31.800 44.800 32.800 45.200 ;
        RECT 33.400 45.100 33.800 45.200 ;
        RECT 33.100 44.800 33.800 45.100 ;
        RECT 27.400 43.800 27.800 44.200 ;
        RECT 29.900 41.100 30.300 44.700 ;
        RECT 32.300 41.100 32.700 44.800 ;
        RECT 33.100 44.200 33.400 44.800 ;
        RECT 33.000 43.800 33.400 44.200 ;
        RECT 34.200 41.400 34.600 45.100 ;
        RECT 35.000 41.700 35.400 45.200 ;
        RECT 35.800 44.800 37.800 45.100 ;
        RECT 35.800 41.400 36.200 44.800 ;
        RECT 34.200 41.100 36.200 41.400 ;
        RECT 37.400 41.100 37.800 44.800 ;
        RECT 39.000 41.100 39.400 49.900 ;
        RECT 41.400 48.900 41.800 49.900 ;
        RECT 39.800 46.800 40.200 47.600 ;
        RECT 41.500 47.200 41.800 48.900 ;
        RECT 43.000 47.900 43.400 49.900 ;
        RECT 43.800 48.000 44.200 49.900 ;
        RECT 45.400 48.000 45.800 49.900 ;
        RECT 47.000 48.900 47.400 49.900 ;
        RECT 47.100 48.100 47.400 48.900 ;
        RECT 49.400 48.900 49.800 49.900 ;
        RECT 51.800 48.900 52.200 49.900 ;
        RECT 48.600 48.100 49.000 48.200 ;
        RECT 43.800 47.900 45.800 48.000 ;
        RECT 43.100 47.200 43.400 47.900 ;
        RECT 43.900 47.700 45.700 47.900 ;
        RECT 47.000 47.800 49.000 48.100 ;
        RECT 45.000 47.200 45.400 47.400 ;
        RECT 47.100 47.200 47.400 47.800 ;
        RECT 41.400 46.800 41.800 47.200 ;
        RECT 43.000 46.800 44.300 47.200 ;
        RECT 45.000 46.900 45.800 47.200 ;
        RECT 45.400 46.800 45.800 46.900 ;
        RECT 47.000 46.800 47.400 47.200 ;
        RECT 41.500 45.100 41.800 46.800 ;
        RECT 42.200 46.100 42.600 46.200 ;
        RECT 42.200 45.800 43.300 46.100 ;
        RECT 42.200 45.400 42.600 45.800 ;
        RECT 43.000 45.200 43.300 45.800 ;
        RECT 43.000 45.100 43.400 45.200 ;
        RECT 44.000 45.100 44.300 46.800 ;
        RECT 47.100 45.100 47.400 46.800 ;
        RECT 49.400 47.200 49.700 48.900 ;
        RECT 50.200 48.100 50.600 48.600 ;
        RECT 51.000 48.100 51.400 48.600 ;
        RECT 51.900 48.200 52.200 48.900 ;
        RECT 50.200 47.800 51.400 48.100 ;
        RECT 51.800 47.800 52.200 48.200 ;
        RECT 53.400 47.900 53.800 49.900 ;
        RECT 54.200 48.000 54.600 49.900 ;
        RECT 55.800 48.000 56.200 49.900 ;
        RECT 54.200 47.900 56.200 48.000 ;
        RECT 51.900 47.200 52.200 47.800 ;
        RECT 53.500 47.200 53.800 47.900 ;
        RECT 54.300 47.700 56.100 47.900 ;
        RECT 49.400 46.800 49.800 47.200 ;
        RECT 51.800 46.800 52.200 47.200 ;
        RECT 53.400 46.800 54.700 47.200 ;
        RECT 49.400 46.200 49.700 46.800 ;
        RECT 47.800 46.100 48.200 46.200 ;
        RECT 48.600 46.100 49.000 46.200 ;
        RECT 47.800 45.800 49.000 46.100 ;
        RECT 47.800 45.400 48.200 45.800 ;
        RECT 48.600 45.400 49.000 45.800 ;
        RECT 49.400 45.800 49.800 46.200 ;
        RECT 49.400 45.100 49.700 45.800 ;
        RECT 51.900 45.100 52.200 46.800 ;
        RECT 54.400 46.200 54.700 46.800 ;
        RECT 52.600 45.400 53.000 46.200 ;
        RECT 54.200 45.800 54.700 46.200 ;
        RECT 53.400 45.100 53.800 45.200 ;
        RECT 54.400 45.100 54.700 45.800 ;
        RECT 41.400 44.700 42.300 45.100 ;
        RECT 43.000 44.800 43.700 45.100 ;
        RECT 44.000 44.800 44.500 45.100 ;
        RECT 41.900 43.200 42.300 44.700 ;
        RECT 43.400 44.200 43.700 44.800 ;
        RECT 43.400 43.800 43.800 44.200 ;
        RECT 41.400 42.800 42.300 43.200 ;
        RECT 41.900 41.100 42.300 42.800 ;
        RECT 44.100 41.100 44.500 44.800 ;
        RECT 47.000 44.700 47.900 45.100 ;
        RECT 47.500 42.200 47.900 44.700 ;
        RECT 48.900 44.700 49.800 45.100 ;
        RECT 51.800 44.700 52.700 45.100 ;
        RECT 53.400 44.800 54.100 45.100 ;
        RECT 54.400 44.800 54.900 45.100 ;
        RECT 47.500 41.800 48.200 42.200 ;
        RECT 47.500 41.100 47.900 41.800 ;
        RECT 48.900 41.100 49.300 44.700 ;
        RECT 52.300 41.100 52.700 44.700 ;
        RECT 53.800 44.200 54.100 44.800 ;
        RECT 53.800 43.800 54.200 44.200 ;
        RECT 54.500 41.100 54.900 44.800 ;
        RECT 56.600 41.100 57.000 49.900 ;
        RECT 58.500 48.200 58.900 49.900 ;
        RECT 63.500 49.200 63.900 49.900 ;
        RECT 63.500 48.800 64.200 49.200 ;
        RECT 63.500 48.200 63.900 48.800 ;
        RECT 58.500 47.900 59.400 48.200 ;
        RECT 57.400 46.800 57.800 47.600 ;
        RECT 59.000 44.100 59.400 47.900 ;
        RECT 63.000 47.900 63.900 48.200 ;
        RECT 65.900 47.900 66.700 49.900 ;
        RECT 62.200 44.100 62.600 44.200 ;
        RECT 59.000 43.800 62.600 44.100 ;
        RECT 59.000 41.100 59.400 43.800 ;
        RECT 63.000 41.100 63.400 47.900 ;
        RECT 65.400 46.800 65.800 47.200 ;
        RECT 65.500 46.600 65.800 46.800 ;
        RECT 65.500 46.200 65.900 46.600 ;
        RECT 66.200 46.200 66.500 47.900 ;
        RECT 66.200 45.800 66.600 46.200 ;
        RECT 67.800 46.100 68.200 46.200 ;
        RECT 67.400 45.800 68.200 46.100 ;
        RECT 66.200 45.700 66.500 45.800 ;
        RECT 65.500 45.400 66.500 45.700 ;
        RECT 67.400 45.600 67.800 45.800 ;
        RECT 63.800 44.400 64.200 45.200 ;
        RECT 65.500 45.100 65.800 45.400 ;
        RECT 64.600 41.400 65.000 45.100 ;
        RECT 65.400 41.700 65.800 45.100 ;
        RECT 66.200 44.800 68.200 45.100 ;
        RECT 66.200 41.400 66.600 44.800 ;
        RECT 64.600 41.100 66.600 41.400 ;
        RECT 67.800 41.100 68.200 44.800 ;
        RECT 69.400 41.100 69.800 49.900 ;
        RECT 71.300 48.200 71.700 49.900 ;
        RECT 71.300 47.900 72.200 48.200 ;
        RECT 70.200 46.800 70.600 47.600 ;
        RECT 71.000 44.400 71.400 45.200 ;
        RECT 71.800 45.100 72.200 47.900 ;
        RECT 72.600 46.800 73.000 47.600 ;
        RECT 74.000 47.100 74.400 49.900 ;
        RECT 77.200 48.200 77.600 49.900 ;
        RECT 81.100 49.200 81.500 49.900 ;
        RECT 81.100 48.800 81.800 49.200 ;
        RECT 81.100 48.200 81.500 48.800 ;
        RECT 82.300 48.200 82.700 48.600 ;
        RECT 77.200 47.800 77.800 48.200 ;
        RECT 80.600 47.900 81.500 48.200 ;
        RECT 77.200 47.100 77.600 47.800 ;
        RECT 73.500 46.900 74.400 47.100 ;
        RECT 76.700 46.900 77.600 47.100 ;
        RECT 73.500 46.800 74.300 46.900 ;
        RECT 76.700 46.800 77.500 46.900 ;
        RECT 79.800 46.800 80.200 47.600 ;
        RECT 72.600 45.800 73.000 46.200 ;
        RECT 72.600 45.100 72.900 45.800 ;
        RECT 73.500 45.200 73.800 46.800 ;
        RECT 74.600 45.800 75.400 46.200 ;
        RECT 71.800 44.800 72.900 45.100 ;
        RECT 73.400 44.800 73.800 45.200 ;
        RECT 75.800 44.800 76.200 45.600 ;
        RECT 76.700 45.200 77.000 46.800 ;
        RECT 77.800 45.800 78.600 46.200 ;
        RECT 76.600 44.800 77.000 45.200 ;
        RECT 79.000 44.800 79.400 45.600 ;
        RECT 71.800 41.100 72.200 44.800 ;
        RECT 73.500 43.500 73.800 44.800 ;
        RECT 74.200 43.800 74.600 44.600 ;
        RECT 76.700 43.500 77.000 44.800 ;
        RECT 77.400 43.800 77.800 44.600 ;
        RECT 73.500 43.200 75.300 43.500 ;
        RECT 76.700 43.200 78.500 43.500 ;
        RECT 73.500 43.100 73.800 43.200 ;
        RECT 73.400 41.100 73.800 43.100 ;
        RECT 75.000 41.100 75.400 43.200 ;
        RECT 76.700 43.100 77.000 43.200 ;
        RECT 76.600 41.100 77.000 43.100 ;
        RECT 78.200 43.100 78.500 43.200 ;
        RECT 78.200 41.100 78.600 43.100 ;
        RECT 80.600 41.100 81.000 47.900 ;
        RECT 82.200 47.800 82.600 48.200 ;
        RECT 83.000 47.900 83.400 49.900 ;
        RECT 85.700 49.200 86.100 49.900 ;
        RECT 85.400 48.800 86.100 49.200 ;
        RECT 85.700 48.200 86.100 48.800 ;
        RECT 85.700 47.900 86.600 48.200 ;
        RECT 82.200 46.100 82.600 46.200 ;
        RECT 83.100 46.100 83.400 47.900 ;
        RECT 83.800 47.100 84.200 47.200 ;
        RECT 85.400 47.100 85.800 47.200 ;
        RECT 83.800 46.800 85.800 47.100 ;
        RECT 83.800 46.400 84.200 46.800 ;
        RECT 84.600 46.100 85.000 46.200 ;
        RECT 82.200 45.800 83.400 46.100 ;
        RECT 84.200 45.800 85.000 46.100 ;
        RECT 81.400 44.400 81.800 45.200 ;
        RECT 82.300 45.100 82.600 45.800 ;
        RECT 84.200 45.600 84.600 45.800 ;
        RECT 82.200 41.100 82.600 45.100 ;
        RECT 83.000 44.800 85.000 45.100 ;
        RECT 83.000 41.100 83.400 44.800 ;
        RECT 84.600 41.100 85.000 44.800 ;
        RECT 85.400 44.400 85.800 45.200 ;
        RECT 86.200 41.100 86.600 47.900 ;
        RECT 87.000 46.800 87.400 47.600 ;
        RECT 0.600 36.200 1.000 39.900 ;
        RECT 1.300 36.200 1.700 36.300 ;
        RECT 0.600 35.900 1.700 36.200 ;
        RECT 2.800 36.200 3.600 39.900 ;
        RECT 4.600 36.200 5.000 36.300 ;
        RECT 5.400 36.200 5.800 39.900 ;
        RECT 6.600 36.800 7.000 37.200 ;
        RECT 6.600 36.200 6.900 36.800 ;
        RECT 7.300 36.200 7.700 39.900 ;
        RECT 2.800 35.900 3.800 36.200 ;
        RECT 4.600 35.900 5.800 36.200 ;
        RECT 6.200 35.900 6.900 36.200 ;
        RECT 7.200 35.900 7.700 36.200 ;
        RECT 1.400 35.600 1.700 35.900 ;
        RECT 1.400 35.300 3.100 35.600 ;
        RECT 2.700 35.200 3.100 35.300 ;
        RECT 3.500 35.200 3.800 35.900 ;
        RECT 6.200 35.800 6.600 35.900 ;
        RECT 3.500 35.100 4.200 35.200 ;
        RECT 6.200 35.100 6.600 35.200 ;
        RECT 1.600 34.900 2.000 35.000 ;
        RECT 3.500 34.900 6.600 35.100 ;
        RECT 1.600 34.600 2.900 34.900 ;
        RECT 2.600 34.300 2.900 34.600 ;
        RECT 3.300 34.800 6.600 34.900 ;
        RECT 3.300 34.600 3.800 34.800 ;
        RECT 2.600 33.900 3.000 34.300 ;
        RECT 1.300 33.400 1.700 33.500 ;
        RECT 0.600 33.100 1.700 33.400 ;
        RECT 0.600 31.100 1.000 33.100 ;
        RECT 3.300 32.900 3.600 34.600 ;
        RECT 7.200 34.200 7.500 35.900 ;
        RECT 7.800 34.400 8.200 35.200 ;
        RECT 6.200 33.800 7.500 34.200 ;
        RECT 8.600 34.100 9.000 34.200 ;
        RECT 8.200 33.800 9.000 34.100 ;
        RECT 4.600 33.400 5.000 33.500 ;
        RECT 4.600 33.100 5.800 33.400 ;
        RECT 6.300 33.100 6.600 33.800 ;
        RECT 8.200 33.600 8.600 33.800 ;
        RECT 9.400 33.400 9.800 34.200 ;
        RECT 7.100 33.100 8.900 33.300 ;
        RECT 10.200 33.100 10.600 39.900 ;
        RECT 11.000 35.800 11.400 36.600 ;
        RECT 13.100 36.200 13.500 39.900 ;
        RECT 13.800 36.800 14.200 37.200 ;
        RECT 13.900 36.200 14.200 36.800 ;
        RECT 16.300 36.300 16.700 39.900 ;
        RECT 13.100 35.900 13.600 36.200 ;
        RECT 13.900 35.900 14.600 36.200 ;
        RECT 15.800 35.900 16.700 36.300 ;
        RECT 18.700 36.200 19.100 39.900 ;
        RECT 19.400 36.800 19.800 37.200 ;
        RECT 19.500 36.200 19.800 36.800 ;
        RECT 20.600 36.200 21.000 39.900 ;
        RECT 22.200 36.200 22.600 39.900 ;
        RECT 18.700 35.900 19.200 36.200 ;
        RECT 19.500 35.900 20.200 36.200 ;
        RECT 20.600 35.900 22.600 36.200 ;
        RECT 23.000 35.900 23.400 39.900 ;
        RECT 24.600 36.100 25.000 36.200 ;
        RECT 25.400 36.100 25.800 39.900 ;
        RECT 11.800 35.100 12.200 35.200 ;
        RECT 12.600 35.100 13.000 35.200 ;
        RECT 11.800 34.800 13.000 35.100 ;
        RECT 12.600 34.400 13.000 34.800 ;
        RECT 13.300 34.200 13.600 35.900 ;
        RECT 14.200 35.800 14.600 35.900 ;
        RECT 14.200 35.100 14.500 35.800 ;
        RECT 15.900 35.100 16.200 35.900 ;
        RECT 14.200 34.800 16.200 35.100 ;
        RECT 16.600 35.100 17.000 35.600 ;
        RECT 18.200 35.100 18.600 35.200 ;
        RECT 16.600 34.800 18.600 35.100 ;
        RECT 15.900 34.200 16.200 34.800 ;
        RECT 18.200 34.400 18.600 34.800 ;
        RECT 18.900 34.200 19.200 35.900 ;
        RECT 19.800 35.800 20.200 35.900 ;
        RECT 21.000 35.200 21.400 35.400 ;
        RECT 23.000 35.200 23.300 35.900 ;
        RECT 24.600 35.800 25.800 36.100 ;
        RECT 20.600 34.900 21.400 35.200 ;
        RECT 22.200 34.900 23.400 35.200 ;
        RECT 20.600 34.800 21.000 34.900 ;
        RECT 11.800 34.100 12.200 34.200 ;
        RECT 11.800 33.800 12.600 34.100 ;
        RECT 13.300 33.800 14.600 34.200 ;
        RECT 15.800 33.800 16.200 34.200 ;
        RECT 17.400 34.100 17.800 34.200 ;
        RECT 17.400 33.800 18.200 34.100 ;
        RECT 18.900 33.800 20.200 34.200 ;
        RECT 20.600 34.100 21.000 34.200 ;
        RECT 21.400 34.100 21.800 34.600 ;
        RECT 20.600 33.800 21.800 34.100 ;
        RECT 12.200 33.600 12.600 33.800 ;
        RECT 11.900 33.100 13.700 33.300 ;
        RECT 14.200 33.100 14.500 33.800 ;
        RECT 2.800 31.100 3.600 32.900 ;
        RECT 5.400 31.100 5.800 33.100 ;
        RECT 6.200 31.100 6.600 33.100 ;
        RECT 7.000 33.000 9.000 33.100 ;
        RECT 7.000 31.100 7.400 33.000 ;
        RECT 8.600 31.100 9.000 33.000 ;
        RECT 10.200 32.800 11.100 33.100 ;
        RECT 10.700 32.200 11.100 32.800 ;
        RECT 11.800 33.000 13.800 33.100 ;
        RECT 10.700 31.800 11.400 32.200 ;
        RECT 10.700 31.100 11.100 31.800 ;
        RECT 11.800 31.100 12.200 33.000 ;
        RECT 13.400 31.100 13.800 33.000 ;
        RECT 14.200 31.100 14.600 33.100 ;
        RECT 15.000 32.400 15.400 33.200 ;
        RECT 15.900 32.100 16.200 33.800 ;
        RECT 17.800 33.600 18.200 33.800 ;
        RECT 17.500 33.100 19.300 33.300 ;
        RECT 19.800 33.100 20.100 33.800 ;
        RECT 22.200 33.100 22.500 34.900 ;
        RECT 23.000 34.800 23.400 34.900 ;
        RECT 15.800 31.100 16.200 32.100 ;
        RECT 17.400 33.000 19.400 33.100 ;
        RECT 17.400 31.100 17.800 33.000 ;
        RECT 19.000 31.100 19.400 33.000 ;
        RECT 19.800 31.100 20.200 33.100 ;
        RECT 22.200 31.100 22.600 33.100 ;
        RECT 23.000 32.800 23.400 33.200 ;
        RECT 22.900 32.400 23.300 32.800 ;
        RECT 25.400 31.100 25.800 35.800 ;
        RECT 27.800 35.100 28.200 39.900 ;
        RECT 28.900 36.300 29.300 39.900 ;
        RECT 28.900 35.900 29.800 36.300 ;
        RECT 28.600 35.100 29.000 35.600 ;
        RECT 27.800 34.800 29.000 35.100 ;
        RECT 26.200 32.400 26.600 33.200 ;
        RECT 27.800 31.100 28.200 34.800 ;
        RECT 29.400 34.200 29.700 35.900 ;
        RECT 31.000 35.800 31.400 36.600 ;
        RECT 28.600 33.800 29.000 34.200 ;
        RECT 29.400 33.800 29.800 34.200 ;
        RECT 28.600 33.100 28.900 33.800 ;
        RECT 29.400 33.100 29.700 33.800 ;
        RECT 28.600 32.800 29.700 33.100 ;
        RECT 29.400 32.100 29.700 32.800 ;
        RECT 30.200 32.400 30.600 33.200 ;
        RECT 31.800 33.100 32.200 39.900 ;
        RECT 33.400 39.600 35.400 39.900 ;
        RECT 33.400 35.900 33.800 39.600 ;
        RECT 34.200 35.900 34.600 39.300 ;
        RECT 35.000 36.200 35.400 39.600 ;
        RECT 36.600 36.200 37.000 39.900 ;
        RECT 35.000 35.900 37.000 36.200 ;
        RECT 37.400 36.200 37.800 39.900 ;
        RECT 39.000 36.200 39.400 39.900 ;
        RECT 37.400 35.900 39.400 36.200 ;
        RECT 39.800 36.100 40.200 39.900 ;
        RECT 34.300 35.600 34.600 35.900 ;
        RECT 39.800 35.800 40.900 36.100 ;
        RECT 34.300 35.300 35.300 35.600 ;
        RECT 35.000 35.200 35.300 35.300 ;
        RECT 36.200 35.200 36.600 35.400 ;
        RECT 37.800 35.200 38.200 35.400 ;
        RECT 39.800 35.200 40.100 35.800 ;
        RECT 40.600 35.200 40.900 35.800 ;
        RECT 35.000 34.800 35.400 35.200 ;
        RECT 36.200 34.900 37.000 35.200 ;
        RECT 36.600 34.800 37.000 34.900 ;
        RECT 37.400 34.900 38.200 35.200 ;
        RECT 39.000 34.900 40.200 35.200 ;
        RECT 37.400 34.800 37.800 34.900 ;
        RECT 34.300 34.400 34.700 34.800 ;
        RECT 34.300 34.200 34.600 34.400 ;
        RECT 34.200 33.800 34.600 34.200 ;
        RECT 35.000 33.100 35.300 34.800 ;
        RECT 35.800 34.100 36.200 34.600 ;
        RECT 37.400 34.100 37.700 34.800 ;
        RECT 35.800 33.800 37.700 34.100 ;
        RECT 38.200 33.800 38.600 34.600 ;
        RECT 39.000 33.100 39.300 34.900 ;
        RECT 39.800 34.800 40.200 34.900 ;
        RECT 40.600 34.800 41.000 35.200 ;
        RECT 41.400 35.100 41.800 39.900 ;
        RECT 42.200 35.800 42.600 36.600 ;
        RECT 44.300 36.200 44.700 39.900 ;
        RECT 45.000 36.800 45.400 37.200 ;
        RECT 45.100 36.200 45.400 36.800 ;
        RECT 46.200 36.200 46.600 39.900 ;
        RECT 47.800 36.200 48.200 39.900 ;
        RECT 44.300 35.900 44.800 36.200 ;
        RECT 45.100 35.900 45.800 36.200 ;
        RECT 46.200 35.900 48.200 36.200 ;
        RECT 48.600 35.900 49.000 39.900 ;
        RECT 43.800 35.100 44.200 35.200 ;
        RECT 41.400 34.800 44.200 35.100 ;
        RECT 40.600 33.400 41.000 34.200 ;
        RECT 31.300 32.800 32.200 33.100 ;
        RECT 31.300 32.200 31.700 32.800 ;
        RECT 34.700 32.200 35.500 33.100 ;
        RECT 29.400 31.100 29.800 32.100 ;
        RECT 31.300 31.800 32.200 32.200 ;
        RECT 34.200 31.800 35.500 32.200 ;
        RECT 31.300 31.100 31.700 31.800 ;
        RECT 34.700 31.100 35.500 31.800 ;
        RECT 39.000 31.100 39.400 33.100 ;
        RECT 39.800 32.800 40.200 33.200 ;
        RECT 41.400 33.100 41.800 34.800 ;
        RECT 43.800 34.400 44.200 34.800 ;
        RECT 44.500 34.200 44.800 35.900 ;
        RECT 45.400 35.800 45.800 35.900 ;
        RECT 45.400 35.100 45.700 35.800 ;
        RECT 46.600 35.200 47.000 35.400 ;
        RECT 48.600 35.200 48.900 35.900 ;
        RECT 46.200 35.100 47.000 35.200 ;
        RECT 45.400 34.900 47.000 35.100 ;
        RECT 47.800 34.900 49.000 35.200 ;
        RECT 45.400 34.800 46.600 34.900 ;
        RECT 43.000 34.100 43.400 34.200 ;
        RECT 43.000 33.800 43.800 34.100 ;
        RECT 44.500 33.800 45.800 34.200 ;
        RECT 47.000 33.800 47.400 34.600 ;
        RECT 43.400 33.600 43.800 33.800 ;
        RECT 43.100 33.100 44.900 33.300 ;
        RECT 45.400 33.200 45.700 33.800 ;
        RECT 41.400 32.800 42.300 33.100 ;
        RECT 39.700 32.400 40.100 32.800 ;
        RECT 41.900 31.100 42.300 32.800 ;
        RECT 43.000 33.000 45.000 33.100 ;
        RECT 43.000 31.100 43.400 33.000 ;
        RECT 44.600 31.100 45.000 33.000 ;
        RECT 45.400 31.100 45.800 33.200 ;
        RECT 47.800 33.100 48.100 34.900 ;
        RECT 48.600 34.800 49.000 34.900 ;
        RECT 48.600 34.200 48.900 34.800 ;
        RECT 48.600 33.800 49.000 34.200 ;
        RECT 48.600 33.100 49.000 33.200 ;
        RECT 49.400 33.100 49.800 39.900 ;
        RECT 51.000 36.200 51.400 39.900 ;
        RECT 52.600 36.200 53.000 39.900 ;
        RECT 51.000 35.900 53.000 36.200 ;
        RECT 53.400 35.900 53.800 39.900 ;
        RECT 55.300 37.200 55.700 39.900 ;
        RECT 54.600 36.800 55.000 37.200 ;
        RECT 55.300 36.800 56.200 37.200 ;
        RECT 54.600 36.200 54.900 36.800 ;
        RECT 55.300 36.200 55.700 36.800 ;
        RECT 54.200 35.900 54.900 36.200 ;
        RECT 55.200 35.900 55.700 36.200 ;
        RECT 51.400 35.200 51.800 35.400 ;
        RECT 53.400 35.200 53.700 35.900 ;
        RECT 54.200 35.800 54.600 35.900 ;
        RECT 50.200 35.100 50.600 35.200 ;
        RECT 51.000 35.100 51.800 35.200 ;
        RECT 50.200 34.900 51.800 35.100 ;
        RECT 52.600 35.100 53.800 35.200 ;
        RECT 54.200 35.100 54.600 35.200 ;
        RECT 52.600 34.900 54.600 35.100 ;
        RECT 50.200 34.800 51.400 34.900 ;
        RECT 51.800 33.800 52.200 34.600 ;
        RECT 47.800 31.100 48.200 33.100 ;
        RECT 48.600 32.800 49.800 33.100 ;
        RECT 48.500 32.400 48.900 32.800 ;
        RECT 49.400 31.100 49.800 32.800 ;
        RECT 50.200 32.400 50.600 33.200 ;
        RECT 52.600 33.100 52.900 34.900 ;
        RECT 53.400 34.800 54.600 34.900 ;
        RECT 55.200 34.200 55.500 35.900 ;
        RECT 55.800 34.400 56.200 35.200 ;
        RECT 54.200 33.800 55.500 34.200 ;
        RECT 56.600 34.100 57.000 34.200 ;
        RECT 56.200 33.800 57.000 34.100 ;
        RECT 52.600 31.100 53.000 33.100 ;
        RECT 53.400 32.800 53.800 33.200 ;
        RECT 54.300 33.100 54.600 33.800 ;
        RECT 56.200 33.600 56.600 33.800 ;
        RECT 57.400 33.400 57.800 34.200 ;
        RECT 55.100 33.100 56.900 33.300 ;
        RECT 53.300 32.400 53.700 32.800 ;
        RECT 54.200 31.100 54.600 33.100 ;
        RECT 55.000 33.000 57.000 33.100 ;
        RECT 55.000 31.100 55.400 33.000 ;
        RECT 56.600 31.100 57.000 33.000 ;
        RECT 58.200 31.100 58.600 39.900 ;
        RECT 60.300 39.200 60.700 39.900 ;
        RECT 59.800 38.800 60.700 39.200 ;
        RECT 60.300 36.200 60.700 38.800 ;
        RECT 61.000 36.800 61.400 37.200 ;
        RECT 61.100 36.200 61.400 36.800 ;
        RECT 65.100 36.200 65.500 39.900 ;
        RECT 65.800 36.800 66.200 37.200 ;
        RECT 65.900 36.200 66.200 36.800 ;
        RECT 67.300 36.300 67.700 39.900 ;
        RECT 60.300 35.900 60.800 36.200 ;
        RECT 61.100 36.100 61.800 36.200 ;
        RECT 63.000 36.100 63.400 36.200 ;
        RECT 61.100 35.900 63.400 36.100 ;
        RECT 65.100 35.900 65.600 36.200 ;
        RECT 65.900 35.900 66.600 36.200 ;
        RECT 67.300 35.900 68.200 36.300 ;
        RECT 70.700 36.200 71.100 39.900 ;
        RECT 71.400 36.800 71.800 37.200 ;
        RECT 71.500 36.200 71.800 36.800 ;
        RECT 70.700 35.900 71.200 36.200 ;
        RECT 71.500 35.900 72.200 36.200 ;
        RECT 59.800 34.400 60.200 35.200 ;
        RECT 60.500 34.200 60.800 35.900 ;
        RECT 61.400 35.800 63.400 35.900 ;
        RECT 64.600 34.400 65.000 35.200 ;
        RECT 65.300 34.200 65.600 35.900 ;
        RECT 66.200 35.800 66.600 35.900 ;
        RECT 67.000 34.800 67.400 35.600 ;
        RECT 67.800 35.100 68.100 35.900 ;
        RECT 70.900 35.200 71.200 35.900 ;
        RECT 71.800 35.800 72.200 35.900 ;
        RECT 68.600 35.100 69.000 35.200 ;
        RECT 67.800 34.800 69.000 35.100 ;
        RECT 69.400 35.100 69.800 35.200 ;
        RECT 70.200 35.100 70.600 35.200 ;
        RECT 69.400 34.800 70.600 35.100 ;
        RECT 67.800 34.200 68.100 34.800 ;
        RECT 70.200 34.400 70.600 34.800 ;
        RECT 70.900 34.800 71.400 35.200 ;
        RECT 73.400 35.100 73.800 39.900 ;
        RECT 75.000 37.900 75.400 39.900 ;
        RECT 75.100 37.800 75.400 37.900 ;
        RECT 76.600 37.900 77.000 39.900 ;
        RECT 79.000 37.900 79.400 39.900 ;
        RECT 76.600 37.800 76.900 37.900 ;
        RECT 75.100 37.500 76.900 37.800 ;
        RECT 79.100 37.800 79.400 37.900 ;
        RECT 80.600 37.900 81.000 39.900 ;
        RECT 80.600 37.800 80.900 37.900 ;
        RECT 79.100 37.500 80.900 37.800 ;
        RECT 74.200 35.800 74.600 36.600 ;
        RECT 75.100 36.200 75.400 37.500 ;
        RECT 75.800 36.400 76.200 37.200 ;
        RECT 76.600 37.100 76.900 37.500 ;
        RECT 76.600 36.800 78.500 37.100 ;
        RECT 78.200 36.200 78.500 36.800 ;
        RECT 79.800 36.400 80.200 37.200 ;
        RECT 80.600 36.200 80.900 37.500 ;
        RECT 82.700 37.200 83.100 39.900 ;
        RECT 82.200 36.800 83.100 37.200 ;
        RECT 83.400 36.800 83.800 37.200 ;
        RECT 82.700 36.200 83.100 36.800 ;
        RECT 83.500 36.200 83.800 36.800 ;
        RECT 84.600 36.200 85.000 39.900 ;
        RECT 75.000 35.800 75.400 36.200 ;
        RECT 73.400 34.800 74.500 35.100 ;
        RECT 70.900 34.200 71.200 34.800 ;
        RECT 59.000 34.100 59.400 34.200 ;
        RECT 59.000 33.800 59.800 34.100 ;
        RECT 60.500 33.800 61.800 34.200 ;
        RECT 62.200 34.100 62.600 34.200 ;
        RECT 63.800 34.100 64.200 34.200 ;
        RECT 62.200 33.800 64.600 34.100 ;
        RECT 65.300 33.800 66.600 34.200 ;
        RECT 67.000 33.800 67.400 34.200 ;
        RECT 67.800 33.800 68.200 34.200 ;
        RECT 68.600 34.100 69.000 34.200 ;
        RECT 69.400 34.100 69.800 34.200 ;
        RECT 68.600 33.800 70.200 34.100 ;
        RECT 70.900 33.800 72.200 34.200 ;
        RECT 59.400 33.600 59.800 33.800 ;
        RECT 59.100 33.100 60.900 33.300 ;
        RECT 61.400 33.100 61.700 33.800 ;
        RECT 64.200 33.600 64.600 33.800 ;
        RECT 63.900 33.100 65.700 33.300 ;
        RECT 66.200 33.100 66.500 33.800 ;
        RECT 67.000 33.100 67.300 33.800 ;
        RECT 59.000 33.000 61.000 33.100 ;
        RECT 59.000 31.100 59.400 33.000 ;
        RECT 60.600 31.100 61.000 33.000 ;
        RECT 61.400 31.100 61.800 33.100 ;
        RECT 63.800 33.000 65.800 33.100 ;
        RECT 63.800 31.100 64.200 33.000 ;
        RECT 65.400 31.100 65.800 33.000 ;
        RECT 66.200 32.800 67.300 33.100 ;
        RECT 66.200 31.100 66.600 32.800 ;
        RECT 67.800 32.100 68.100 33.800 ;
        RECT 69.800 33.600 70.200 33.800 ;
        RECT 68.600 32.400 69.000 33.200 ;
        RECT 69.500 33.100 71.300 33.300 ;
        RECT 71.800 33.100 72.100 33.800 ;
        RECT 72.600 33.400 73.000 34.200 ;
        RECT 73.400 33.100 73.800 34.800 ;
        RECT 74.200 34.200 74.500 34.800 ;
        RECT 75.100 34.200 75.400 35.800 ;
        RECT 77.400 35.400 77.800 36.200 ;
        RECT 78.200 35.400 78.600 36.200 ;
        RECT 80.600 35.800 81.000 36.200 ;
        RECT 82.700 35.900 83.200 36.200 ;
        RECT 83.500 35.900 84.200 36.200 ;
        RECT 84.600 35.900 85.700 36.200 ;
        RECT 76.200 34.800 77.000 35.200 ;
        RECT 79.000 34.800 79.800 35.200 ;
        RECT 80.600 34.200 80.900 35.800 ;
        RECT 82.200 34.400 82.600 35.200 ;
        RECT 82.900 34.200 83.200 35.900 ;
        RECT 83.800 35.800 84.200 35.900 ;
        RECT 85.400 35.600 85.700 35.900 ;
        RECT 85.400 35.200 86.000 35.600 ;
        RECT 84.600 34.400 85.000 35.200 ;
        RECT 74.200 33.800 74.600 34.200 ;
        RECT 75.100 34.100 75.900 34.200 ;
        RECT 80.100 34.100 81.000 34.200 ;
        RECT 75.100 33.900 76.000 34.100 ;
        RECT 69.400 33.000 71.400 33.100 ;
        RECT 67.800 31.100 68.200 32.100 ;
        RECT 69.400 31.100 69.800 33.000 ;
        RECT 71.000 31.100 71.400 33.000 ;
        RECT 71.800 31.100 72.200 33.100 ;
        RECT 73.400 32.800 74.300 33.100 ;
        RECT 73.900 31.100 74.300 32.800 ;
        RECT 75.600 31.100 76.000 33.900 ;
        RECT 80.000 33.800 81.000 34.100 ;
        RECT 81.400 34.100 81.800 34.200 ;
        RECT 81.400 33.800 82.200 34.100 ;
        RECT 82.900 33.800 84.200 34.200 ;
        RECT 80.000 31.100 80.400 33.800 ;
        RECT 81.800 33.600 82.200 33.800 ;
        RECT 81.500 33.100 83.300 33.300 ;
        RECT 83.800 33.100 84.100 33.800 ;
        RECT 85.400 33.700 85.700 35.200 ;
        RECT 84.600 33.400 85.700 33.700 ;
        RECT 81.400 33.000 83.400 33.100 ;
        RECT 81.400 31.100 81.800 33.000 ;
        RECT 83.000 31.100 83.400 33.000 ;
        RECT 83.800 31.100 84.200 33.100 ;
        RECT 84.600 31.100 85.000 33.400 ;
        RECT 0.600 27.900 1.000 29.900 ;
        RECT 2.800 28.100 3.600 29.900 ;
        RECT 0.600 27.600 1.900 27.900 ;
        RECT 1.500 27.500 1.900 27.600 ;
        RECT 2.200 27.400 3.000 27.800 ;
        RECT 3.300 27.100 3.600 28.100 ;
        RECT 5.400 27.900 5.800 29.900 ;
        RECT 6.500 29.200 6.900 29.900 ;
        RECT 6.500 28.800 7.400 29.200 ;
        RECT 6.500 28.200 6.900 28.800 ;
        RECT 6.500 27.900 7.400 28.200 ;
        RECT 3.900 27.400 4.300 27.800 ;
        RECT 4.600 27.600 5.800 27.900 ;
        RECT 4.600 27.500 5.000 27.600 ;
        RECT 3.100 26.800 3.600 27.100 ;
        RECT 4.000 27.200 4.300 27.400 ;
        RECT 4.000 26.800 4.400 27.200 ;
        RECT 3.100 26.200 3.400 26.800 ;
        RECT 1.700 26.100 2.100 26.200 ;
        RECT 1.700 25.800 2.500 26.100 ;
        RECT 3.000 25.800 3.400 26.200 ;
        RECT 2.100 25.700 2.500 25.800 ;
        RECT 3.100 25.100 3.400 25.800 ;
        RECT 0.600 24.800 1.900 25.100 ;
        RECT 0.600 21.100 1.000 24.800 ;
        RECT 1.500 24.700 1.900 24.800 ;
        RECT 2.800 22.200 3.600 25.100 ;
        RECT 4.600 24.800 5.800 25.100 ;
        RECT 4.600 24.700 5.000 24.800 ;
        RECT 2.800 21.800 4.200 22.200 ;
        RECT 2.800 21.100 3.600 21.800 ;
        RECT 5.400 21.100 5.800 24.800 ;
        RECT 6.200 24.400 6.600 25.200 ;
        RECT 7.000 21.100 7.400 27.900 ;
        RECT 7.800 26.800 8.200 27.600 ;
        RECT 10.400 27.100 10.800 29.900 ;
        RECT 11.800 28.000 12.200 29.900 ;
        RECT 13.400 28.000 13.800 29.900 ;
        RECT 11.800 27.900 13.800 28.000 ;
        RECT 14.200 27.900 14.600 29.900 ;
        RECT 15.800 28.900 16.200 29.900 ;
        RECT 11.900 27.700 13.700 27.900 ;
        RECT 12.200 27.200 12.600 27.400 ;
        RECT 14.200 27.200 14.500 27.900 ;
        RECT 15.000 27.800 15.400 28.600 ;
        RECT 15.900 27.200 16.200 28.900 ;
        RECT 17.400 28.000 17.800 29.900 ;
        RECT 19.000 28.000 19.400 29.900 ;
        RECT 17.400 27.900 19.400 28.000 ;
        RECT 19.800 27.900 20.200 29.900 ;
        RECT 20.600 28.000 21.000 29.900 ;
        RECT 22.200 28.000 22.600 29.900 ;
        RECT 20.600 27.900 22.600 28.000 ;
        RECT 23.000 27.900 23.400 29.900 ;
        RECT 25.400 27.900 25.800 29.900 ;
        RECT 26.200 28.000 26.600 29.900 ;
        RECT 27.800 28.000 28.200 29.900 ;
        RECT 29.400 28.900 29.800 29.900 ;
        RECT 26.200 27.900 28.200 28.000 ;
        RECT 17.500 27.700 19.300 27.900 ;
        RECT 17.800 27.200 18.200 27.400 ;
        RECT 19.800 27.200 20.100 27.900 ;
        RECT 20.700 27.700 22.500 27.900 ;
        RECT 21.000 27.200 21.400 27.400 ;
        RECT 23.000 27.200 23.300 27.900 ;
        RECT 25.500 27.200 25.800 27.900 ;
        RECT 26.300 27.700 28.100 27.900 ;
        RECT 29.500 27.200 29.800 28.900 ;
        RECT 30.200 28.100 30.600 28.200 ;
        RECT 31.000 28.100 31.400 29.900 ;
        RECT 30.200 27.800 31.400 28.100 ;
        RECT 32.600 28.000 33.000 29.900 ;
        RECT 34.200 28.000 34.600 29.900 ;
        RECT 32.600 27.900 34.600 28.000 ;
        RECT 35.000 27.900 35.400 29.900 ;
        RECT 37.100 27.900 37.900 29.900 ;
        RECT 40.600 28.900 41.000 29.900 ;
        RECT 10.400 26.900 11.300 27.100 ;
        RECT 10.500 26.800 11.300 26.900 ;
        RECT 11.800 26.900 12.600 27.200 ;
        RECT 11.800 26.800 12.200 26.900 ;
        RECT 13.300 26.800 14.600 27.200 ;
        RECT 15.800 27.100 16.200 27.200 ;
        RECT 17.400 27.100 18.200 27.200 ;
        RECT 15.800 26.900 18.200 27.100 ;
        RECT 15.800 26.800 17.800 26.900 ;
        RECT 18.900 26.800 20.200 27.200 ;
        RECT 20.600 26.900 21.400 27.200 ;
        RECT 20.600 26.800 21.000 26.900 ;
        RECT 22.100 26.800 23.400 27.200 ;
        RECT 25.400 26.800 26.700 27.200 ;
        RECT 29.400 26.800 29.800 27.200 ;
        RECT 9.400 25.800 10.600 26.200 ;
        RECT 8.600 24.800 9.000 25.600 ;
        RECT 11.000 25.200 11.300 26.800 ;
        RECT 12.600 25.800 13.000 26.600 ;
        RECT 13.300 26.100 13.600 26.800 ;
        RECT 15.000 26.100 15.400 26.200 ;
        RECT 13.300 25.800 15.400 26.100 ;
        RECT 11.000 24.800 11.400 25.200 ;
        RECT 13.300 25.100 13.600 25.800 ;
        RECT 14.200 25.100 14.600 25.200 ;
        RECT 15.900 25.100 16.200 26.800 ;
        RECT 16.600 25.400 17.000 26.200 ;
        RECT 18.200 25.800 18.600 26.600 ;
        RECT 18.900 25.100 19.200 26.800 ;
        RECT 21.400 25.800 21.800 26.600 ;
        RECT 19.800 25.100 20.200 25.200 ;
        RECT 22.100 25.100 22.400 26.800 ;
        RECT 26.400 26.100 26.700 26.800 ;
        RECT 23.000 25.800 26.700 26.100 ;
        RECT 23.000 25.200 23.300 25.800 ;
        RECT 23.000 25.100 23.400 25.200 ;
        RECT 13.100 24.800 13.600 25.100 ;
        RECT 13.900 24.800 14.600 25.100 ;
        RECT 10.200 23.800 10.600 24.600 ;
        RECT 11.000 23.500 11.300 24.800 ;
        RECT 9.500 23.200 11.300 23.500 ;
        RECT 9.500 23.100 9.800 23.200 ;
        RECT 9.400 21.100 9.800 23.100 ;
        RECT 11.000 23.100 11.300 23.200 ;
        RECT 11.000 21.100 11.400 23.100 ;
        RECT 13.100 21.100 13.500 24.800 ;
        RECT 13.900 24.200 14.200 24.800 ;
        RECT 15.800 24.700 16.700 25.100 ;
        RECT 13.800 23.800 14.200 24.200 ;
        RECT 16.300 21.100 16.700 24.700 ;
        RECT 18.700 24.800 19.200 25.100 ;
        RECT 19.500 24.800 20.200 25.100 ;
        RECT 21.900 24.800 22.400 25.100 ;
        RECT 22.700 24.800 23.400 25.100 ;
        RECT 25.400 25.100 25.800 25.200 ;
        RECT 26.400 25.100 26.700 25.800 ;
        RECT 29.500 25.100 29.800 26.800 ;
        RECT 30.200 26.100 30.600 26.200 ;
        RECT 31.000 26.100 31.400 27.800 ;
        RECT 32.700 27.700 34.500 27.900 ;
        RECT 33.000 27.200 33.400 27.400 ;
        RECT 35.000 27.200 35.300 27.900 ;
        RECT 32.600 26.900 33.400 27.200 ;
        RECT 32.600 26.800 33.000 26.900 ;
        RECT 34.100 26.800 35.400 27.200 ;
        RECT 36.600 26.800 37.000 27.200 ;
        RECT 30.200 25.800 31.400 26.100 ;
        RECT 33.400 25.800 33.800 26.600 ;
        RECT 30.200 25.400 30.600 25.800 ;
        RECT 25.400 24.800 26.100 25.100 ;
        RECT 26.400 24.800 26.900 25.100 ;
        RECT 18.700 22.200 19.100 24.800 ;
        RECT 19.500 24.200 19.800 24.800 ;
        RECT 19.400 23.800 19.800 24.200 ;
        RECT 21.900 22.200 22.300 24.800 ;
        RECT 22.700 24.200 23.000 24.800 ;
        RECT 22.600 23.800 23.000 24.200 ;
        RECT 25.800 24.200 26.100 24.800 ;
        RECT 25.800 23.800 26.200 24.200 ;
        RECT 18.200 21.800 19.100 22.200 ;
        RECT 21.400 21.800 22.300 22.200 ;
        RECT 18.700 21.100 19.100 21.800 ;
        RECT 21.900 21.100 22.300 21.800 ;
        RECT 26.500 21.100 26.900 24.800 ;
        RECT 29.400 24.700 30.300 25.100 ;
        RECT 29.900 22.200 30.300 24.700 ;
        RECT 29.400 21.800 30.300 22.200 ;
        RECT 29.900 21.100 30.300 21.800 ;
        RECT 31.000 21.100 31.400 25.800 ;
        RECT 34.100 25.100 34.400 26.800 ;
        RECT 36.700 26.600 37.000 26.800 ;
        RECT 36.700 26.200 37.100 26.600 ;
        RECT 37.400 26.200 37.700 27.900 ;
        RECT 39.800 27.800 40.200 28.600 ;
        RECT 40.700 27.200 41.000 28.900 ;
        RECT 43.800 27.900 44.200 29.900 ;
        RECT 44.500 28.200 44.900 28.600 ;
        RECT 38.200 26.400 38.600 27.200 ;
        RECT 40.600 27.100 41.000 27.200 ;
        RECT 40.600 26.800 42.500 27.100 ;
        RECT 37.400 25.800 37.800 26.200 ;
        RECT 39.000 26.100 39.400 26.200 ;
        RECT 38.600 25.800 39.400 26.100 ;
        RECT 37.400 25.700 37.700 25.800 ;
        RECT 36.700 25.400 37.700 25.700 ;
        RECT 38.600 25.600 39.000 25.800 ;
        RECT 35.000 25.100 35.400 25.200 ;
        RECT 36.700 25.100 37.000 25.400 ;
        RECT 40.700 25.100 41.000 26.800 ;
        RECT 42.200 26.200 42.500 26.800 ;
        RECT 43.000 26.400 43.400 27.200 ;
        RECT 41.400 25.400 41.800 26.200 ;
        RECT 42.200 26.100 42.600 26.200 ;
        RECT 43.800 26.100 44.100 27.900 ;
        RECT 44.600 27.800 45.000 28.200 ;
        RECT 45.400 28.000 45.800 29.900 ;
        RECT 47.000 28.000 47.400 29.900 ;
        RECT 45.400 27.900 47.400 28.000 ;
        RECT 47.800 27.900 48.200 29.900 ;
        RECT 50.200 27.900 50.600 29.900 ;
        RECT 50.900 28.200 51.300 28.600 ;
        RECT 45.500 27.700 47.300 27.900 ;
        RECT 45.800 27.200 46.200 27.400 ;
        RECT 47.800 27.200 48.100 27.900 ;
        RECT 45.400 26.900 46.200 27.200 ;
        RECT 45.400 26.800 45.800 26.900 ;
        RECT 46.900 26.800 48.200 27.200 ;
        RECT 44.600 26.100 45.000 26.200 ;
        RECT 42.200 25.800 43.000 26.100 ;
        RECT 43.800 25.800 45.000 26.100 ;
        RECT 46.200 25.800 46.600 26.600 ;
        RECT 42.600 25.600 43.000 25.800 ;
        RECT 44.600 25.100 44.900 25.800 ;
        RECT 46.900 25.100 47.200 26.800 ;
        RECT 49.400 26.400 49.800 27.200 ;
        RECT 48.600 26.100 49.000 26.200 ;
        RECT 50.200 26.100 50.500 27.900 ;
        RECT 51.000 27.800 51.400 28.200 ;
        RECT 51.800 27.800 52.200 28.600 ;
        RECT 52.600 27.100 53.000 29.900 ;
        RECT 53.400 29.600 55.400 29.900 ;
        RECT 53.400 27.900 53.800 29.600 ;
        RECT 54.200 27.900 54.600 29.300 ;
        RECT 55.000 28.000 55.400 29.600 ;
        RECT 56.600 28.000 57.000 29.900 ;
        RECT 58.700 28.200 59.100 29.900 ;
        RECT 62.200 28.900 62.600 29.900 ;
        RECT 55.000 27.900 57.000 28.000 ;
        RECT 58.200 27.900 59.100 28.200 ;
        RECT 59.800 28.100 60.200 28.200 ;
        RECT 62.200 28.100 62.500 28.900 ;
        RECT 54.200 27.200 54.500 27.900 ;
        RECT 55.100 27.700 56.900 27.900 ;
        RECT 56.200 27.200 56.600 27.400 ;
        RECT 53.400 27.100 53.800 27.200 ;
        RECT 52.600 26.800 53.800 27.100 ;
        RECT 54.200 26.900 55.400 27.200 ;
        RECT 56.200 26.900 57.000 27.200 ;
        RECT 55.000 26.800 55.400 26.900 ;
        RECT 56.600 26.800 57.000 26.900 ;
        RECT 57.400 26.800 57.800 27.600 ;
        RECT 51.000 26.100 51.400 26.200 ;
        RECT 48.600 25.800 49.400 26.100 ;
        RECT 50.200 25.800 51.400 26.100 ;
        RECT 49.000 25.600 49.400 25.800 ;
        RECT 47.800 25.100 48.200 25.200 ;
        RECT 51.000 25.100 51.300 25.800 ;
        RECT 33.900 24.800 34.400 25.100 ;
        RECT 34.700 24.800 35.400 25.100 ;
        RECT 33.900 21.100 34.300 24.800 ;
        RECT 34.700 24.200 35.000 24.800 ;
        RECT 34.600 23.800 35.000 24.200 ;
        RECT 35.800 21.400 36.200 25.100 ;
        RECT 36.600 21.700 37.000 25.100 ;
        RECT 37.400 24.800 39.400 25.100 ;
        RECT 37.400 21.400 37.800 24.800 ;
        RECT 35.800 21.100 37.800 21.400 ;
        RECT 39.000 21.100 39.400 24.800 ;
        RECT 40.600 24.700 41.500 25.100 ;
        RECT 41.100 21.100 41.500 24.700 ;
        RECT 42.200 24.800 44.200 25.100 ;
        RECT 42.200 21.100 42.600 24.800 ;
        RECT 43.800 21.100 44.200 24.800 ;
        RECT 44.600 21.100 45.000 25.100 ;
        RECT 46.700 24.800 47.200 25.100 ;
        RECT 47.500 24.800 48.200 25.100 ;
        RECT 48.600 24.800 50.600 25.100 ;
        RECT 46.700 22.200 47.100 24.800 ;
        RECT 47.500 24.200 47.800 24.800 ;
        RECT 47.400 23.800 47.800 24.200 ;
        RECT 46.200 21.800 47.100 22.200 ;
        RECT 46.700 21.100 47.100 21.800 ;
        RECT 48.600 21.100 49.000 24.800 ;
        RECT 50.200 21.100 50.600 24.800 ;
        RECT 51.000 24.100 51.400 25.100 ;
        RECT 51.800 24.100 52.200 24.200 ;
        RECT 51.000 23.800 52.200 24.100 ;
        RECT 51.000 21.100 51.400 23.800 ;
        RECT 52.600 21.100 53.000 26.800 ;
        RECT 53.400 26.400 53.800 26.800 ;
        RECT 54.200 25.800 54.600 26.600 ;
        RECT 55.100 25.100 55.400 26.800 ;
        RECT 55.800 26.100 56.200 26.600 ;
        RECT 56.600 26.100 57.000 26.200 ;
        RECT 55.800 25.800 57.000 26.100 ;
        RECT 58.200 26.100 58.600 27.900 ;
        RECT 59.800 27.800 62.500 28.100 ;
        RECT 63.000 27.800 63.400 28.600 ;
        RECT 63.800 28.000 64.200 29.900 ;
        RECT 65.400 28.000 65.800 29.900 ;
        RECT 63.800 27.900 65.800 28.000 ;
        RECT 66.200 27.900 66.600 29.900 ;
        RECT 67.300 28.200 67.700 29.900 ;
        RECT 69.700 28.200 70.100 29.900 ;
        RECT 67.300 27.900 68.200 28.200 ;
        RECT 69.700 27.900 70.600 28.200 ;
        RECT 62.200 27.200 62.500 27.800 ;
        RECT 63.900 27.700 65.700 27.900 ;
        RECT 64.200 27.200 64.600 27.400 ;
        RECT 66.200 27.200 66.500 27.900 ;
        RECT 62.200 26.800 62.600 27.200 ;
        RECT 63.800 26.900 64.600 27.200 ;
        RECT 63.800 26.800 64.200 26.900 ;
        RECT 65.300 26.800 66.600 27.200 ;
        RECT 61.400 26.100 61.800 26.200 ;
        RECT 58.200 25.800 61.800 26.100 ;
        RECT 54.700 22.200 55.700 25.100 ;
        RECT 54.700 21.800 56.200 22.200 ;
        RECT 54.700 21.100 55.700 21.800 ;
        RECT 58.200 21.100 58.600 25.800 ;
        RECT 61.400 25.400 61.800 25.800 ;
        RECT 59.000 24.400 59.400 25.200 ;
        RECT 62.200 25.100 62.500 26.800 ;
        RECT 64.600 25.800 65.000 26.600 ;
        RECT 65.300 25.100 65.600 26.800 ;
        RECT 67.800 26.100 68.200 27.900 ;
        RECT 68.600 27.100 69.000 27.600 ;
        RECT 70.200 27.100 70.600 27.900 ;
        RECT 68.600 26.800 70.600 27.100 ;
        RECT 71.000 26.800 71.400 27.600 ;
        RECT 69.400 26.100 69.800 26.200 ;
        RECT 67.800 25.800 69.800 26.100 ;
        RECT 66.200 25.100 66.600 25.200 ;
        RECT 61.700 24.700 62.600 25.100 ;
        RECT 65.100 24.800 65.600 25.100 ;
        RECT 65.900 24.800 66.600 25.100 ;
        RECT 61.700 21.100 62.100 24.700 ;
        RECT 65.100 21.100 65.500 24.800 ;
        RECT 65.900 24.200 66.200 24.800 ;
        RECT 67.000 24.400 67.400 25.200 ;
        RECT 65.800 23.800 66.200 24.200 ;
        RECT 67.800 21.100 68.200 25.800 ;
        RECT 69.400 24.400 69.800 25.200 ;
        RECT 70.200 21.100 70.600 26.800 ;
        RECT 72.600 21.100 73.000 29.900 ;
        RECT 74.200 27.800 74.600 28.600 ;
        RECT 73.400 26.800 73.800 27.600 ;
        RECT 75.000 26.100 75.400 29.900 ;
        RECT 77.400 27.900 77.800 29.900 ;
        RECT 78.100 28.200 78.500 28.600 ;
        RECT 78.200 28.100 78.600 28.200 ;
        RECT 79.000 28.100 79.400 28.600 ;
        RECT 76.600 26.400 77.000 27.200 ;
        RECT 75.800 26.100 76.200 26.200 ;
        RECT 77.400 26.100 77.700 27.900 ;
        RECT 78.200 27.800 79.400 28.100 ;
        RECT 78.200 26.100 78.600 26.200 ;
        RECT 75.000 25.800 76.600 26.100 ;
        RECT 77.400 25.800 78.600 26.100 ;
        RECT 75.000 21.100 75.400 25.800 ;
        RECT 76.200 25.600 76.600 25.800 ;
        RECT 78.200 25.100 78.500 25.800 ;
        RECT 75.800 24.800 77.800 25.100 ;
        RECT 75.800 21.100 76.200 24.800 ;
        RECT 77.400 21.100 77.800 24.800 ;
        RECT 78.200 21.100 78.600 25.100 ;
        RECT 79.800 21.100 80.200 29.900 ;
        RECT 80.600 28.000 81.000 29.900 ;
        RECT 82.200 28.000 82.600 29.900 ;
        RECT 80.600 27.900 82.600 28.000 ;
        RECT 83.000 27.900 83.400 29.900 ;
        RECT 85.100 28.200 85.500 29.900 ;
        RECT 84.600 27.900 85.500 28.200 ;
        RECT 80.700 27.700 82.500 27.900 ;
        RECT 81.000 27.200 81.400 27.400 ;
        RECT 83.000 27.200 83.300 27.900 ;
        RECT 80.600 26.900 81.400 27.200 ;
        RECT 80.600 26.800 81.000 26.900 ;
        RECT 82.100 26.800 83.400 27.200 ;
        RECT 81.400 25.800 81.800 26.600 ;
        RECT 82.100 25.100 82.400 26.800 ;
        RECT 83.000 25.100 83.400 25.200 ;
        RECT 81.900 24.800 82.400 25.100 ;
        RECT 82.700 24.800 83.400 25.100 ;
        RECT 81.900 21.100 82.300 24.800 ;
        RECT 82.700 24.200 83.000 24.800 ;
        RECT 82.600 23.800 83.000 24.200 ;
        RECT 84.600 21.100 85.000 27.900 ;
        RECT 2.200 16.200 2.600 19.900 ;
        RECT 3.000 17.900 3.400 19.900 ;
        RECT 3.100 17.800 3.400 17.900 ;
        RECT 4.600 17.900 5.000 19.900 ;
        RECT 4.600 17.800 4.900 17.900 ;
        RECT 3.100 17.500 4.900 17.800 ;
        RECT 3.100 16.200 3.400 17.500 ;
        RECT 3.800 16.400 4.200 17.200 ;
        RECT 7.500 16.200 7.900 19.900 ;
        RECT 8.200 16.800 8.600 17.200 ;
        RECT 8.300 16.200 8.600 16.800 ;
        RECT 1.500 15.900 2.600 16.200 ;
        RECT 1.500 15.600 1.800 15.900 ;
        RECT 3.000 15.800 3.400 16.200 ;
        RECT 1.200 15.200 1.800 15.600 ;
        RECT 1.500 13.700 1.800 15.200 ;
        RECT 2.200 15.100 2.600 15.200 ;
        RECT 3.100 15.100 3.400 15.800 ;
        RECT 5.400 15.400 5.800 16.200 ;
        RECT 7.000 15.800 8.000 16.200 ;
        RECT 8.300 16.100 9.000 16.200 ;
        RECT 9.400 16.100 9.800 19.900 ;
        RECT 8.300 15.900 9.800 16.100 ;
        RECT 10.200 16.200 10.600 19.900 ;
        RECT 11.800 16.200 12.200 19.900 ;
        RECT 10.200 15.900 12.200 16.200 ;
        RECT 13.900 16.200 14.300 19.900 ;
        RECT 14.600 16.800 15.000 17.200 ;
        RECT 14.700 16.200 15.000 16.800 ;
        RECT 16.100 16.300 16.500 19.900 ;
        RECT 13.900 15.900 14.400 16.200 ;
        RECT 14.700 15.900 15.400 16.200 ;
        RECT 16.100 15.900 17.000 16.300 ;
        RECT 19.500 16.200 19.900 19.900 ;
        RECT 20.200 16.800 20.600 17.200 ;
        RECT 20.300 16.200 20.600 16.800 ;
        RECT 22.700 16.300 23.100 19.900 ;
        RECT 19.500 15.900 20.000 16.200 ;
        RECT 20.300 15.900 21.000 16.200 ;
        RECT 8.600 15.800 9.800 15.900 ;
        RECT 2.200 14.800 3.400 15.100 ;
        RECT 4.200 14.800 5.000 15.200 ;
        RECT 6.200 15.100 6.600 15.200 ;
        RECT 7.000 15.100 7.400 15.200 ;
        RECT 6.200 14.800 7.400 15.100 ;
        RECT 2.200 14.400 2.600 14.800 ;
        RECT 3.100 14.200 3.400 14.800 ;
        RECT 7.000 14.400 7.400 14.800 ;
        RECT 7.700 14.200 8.000 15.800 ;
        RECT 9.500 15.200 9.800 15.800 ;
        RECT 11.400 15.200 11.800 15.400 ;
        RECT 9.400 14.900 10.600 15.200 ;
        RECT 11.400 15.100 12.200 15.200 ;
        RECT 12.600 15.100 13.000 15.200 ;
        RECT 11.400 14.900 13.000 15.100 ;
        RECT 9.400 14.800 9.800 14.900 ;
        RECT 3.100 14.100 3.900 14.200 ;
        RECT 6.200 14.100 6.600 14.200 ;
        RECT 3.100 13.900 4.000 14.100 ;
        RECT 1.500 13.400 2.600 13.700 ;
        RECT 2.200 11.100 2.600 13.400 ;
        RECT 3.600 11.100 4.000 13.900 ;
        RECT 6.200 13.800 7.000 14.100 ;
        RECT 7.700 13.800 9.000 14.200 ;
        RECT 6.600 13.600 7.000 13.800 ;
        RECT 6.300 13.100 8.100 13.300 ;
        RECT 8.600 13.100 8.900 13.800 ;
        RECT 6.200 13.000 8.200 13.100 ;
        RECT 6.200 11.100 6.600 13.000 ;
        RECT 7.800 11.100 8.200 13.000 ;
        RECT 8.600 11.100 9.000 13.100 ;
        RECT 9.400 12.800 9.800 13.200 ;
        RECT 10.300 13.100 10.600 14.900 ;
        RECT 11.800 14.800 13.000 14.900 ;
        RECT 11.000 13.800 11.400 14.600 ;
        RECT 12.600 14.200 12.900 14.800 ;
        RECT 13.400 14.400 13.800 15.200 ;
        RECT 14.100 14.200 14.400 15.900 ;
        RECT 15.000 15.800 15.400 15.900 ;
        RECT 15.800 14.800 16.200 15.600 ;
        RECT 16.600 14.200 16.900 15.900 ;
        RECT 19.000 14.400 19.400 15.200 ;
        RECT 19.700 14.200 20.000 15.900 ;
        RECT 20.600 15.800 21.000 15.900 ;
        RECT 22.200 15.900 23.100 16.300 ;
        RECT 25.800 16.800 26.200 17.200 ;
        RECT 25.800 16.200 26.100 16.800 ;
        RECT 26.500 16.200 26.900 19.900 ;
        RECT 25.400 15.900 26.100 16.200 ;
        RECT 26.400 15.900 26.900 16.200 ;
        RECT 28.600 16.200 29.000 19.900 ;
        RECT 30.200 16.200 30.600 19.900 ;
        RECT 28.600 15.900 30.600 16.200 ;
        RECT 31.000 15.900 31.400 19.900 ;
        RECT 33.100 16.200 33.500 19.900 ;
        RECT 33.800 16.800 34.200 17.200 ;
        RECT 33.900 16.200 34.200 16.800 ;
        RECT 22.200 15.800 22.600 15.900 ;
        RECT 25.400 15.800 25.800 15.900 ;
        RECT 22.300 14.200 22.600 15.800 ;
        RECT 23.000 14.800 23.400 15.600 ;
        RECT 24.600 15.100 25.000 15.200 ;
        RECT 26.400 15.100 26.700 15.900 ;
        RECT 29.000 15.200 29.400 15.400 ;
        RECT 31.000 15.200 31.300 15.900 ;
        RECT 32.600 15.800 33.600 16.200 ;
        RECT 33.900 15.900 34.600 16.200 ;
        RECT 34.200 15.800 34.600 15.900 ;
        RECT 24.600 14.800 26.700 15.100 ;
        RECT 28.600 14.900 29.400 15.200 ;
        RECT 30.200 14.900 31.400 15.200 ;
        RECT 28.600 14.800 29.000 14.900 ;
        RECT 26.400 14.200 26.700 14.800 ;
        RECT 12.600 14.100 13.000 14.200 ;
        RECT 12.600 13.800 13.400 14.100 ;
        RECT 14.100 13.800 15.400 14.200 ;
        RECT 16.600 13.800 17.000 14.200 ;
        RECT 18.200 14.100 18.600 14.200 ;
        RECT 18.200 13.800 19.000 14.100 ;
        RECT 19.700 13.800 21.000 14.200 ;
        RECT 22.200 13.800 22.600 14.200 ;
        RECT 25.400 13.800 26.700 14.200 ;
        RECT 29.400 13.800 29.800 14.600 ;
        RECT 13.000 13.600 13.400 13.800 ;
        RECT 12.700 13.100 14.500 13.300 ;
        RECT 15.000 13.100 15.300 13.800 ;
        RECT 9.500 12.400 9.900 12.800 ;
        RECT 10.200 11.100 10.600 13.100 ;
        RECT 12.600 13.000 14.600 13.100 ;
        RECT 12.600 11.100 13.000 13.000 ;
        RECT 14.200 11.100 14.600 13.000 ;
        RECT 15.000 11.100 15.400 13.100 ;
        RECT 16.600 12.200 16.900 13.800 ;
        RECT 18.600 13.600 19.000 13.800 ;
        RECT 17.400 12.400 17.800 13.200 ;
        RECT 18.300 13.100 20.100 13.300 ;
        RECT 20.600 13.100 20.900 13.800 ;
        RECT 18.200 13.000 20.200 13.100 ;
        RECT 16.600 11.100 17.000 12.200 ;
        RECT 18.200 11.100 18.600 13.000 ;
        RECT 19.800 11.100 20.200 13.000 ;
        RECT 20.600 11.100 21.000 13.100 ;
        RECT 21.400 12.400 21.800 13.200 ;
        RECT 22.300 12.100 22.600 13.800 ;
        RECT 25.500 13.100 25.800 13.800 ;
        RECT 26.300 13.100 28.100 13.300 ;
        RECT 30.200 13.100 30.500 14.900 ;
        RECT 31.000 14.800 31.400 14.900 ;
        RECT 32.600 14.400 33.000 15.200 ;
        RECT 33.300 14.200 33.600 15.800 ;
        RECT 31.800 14.100 32.200 14.200 ;
        RECT 31.800 13.800 32.600 14.100 ;
        RECT 33.300 13.800 34.600 14.200 ;
        RECT 32.200 13.600 32.600 13.800 ;
        RECT 22.200 11.100 22.600 12.100 ;
        RECT 25.400 11.100 25.800 13.100 ;
        RECT 26.200 13.000 28.200 13.100 ;
        RECT 26.200 11.100 26.600 13.000 ;
        RECT 27.800 11.100 28.200 13.000 ;
        RECT 30.200 11.100 30.600 13.100 ;
        RECT 31.000 12.800 31.400 13.200 ;
        RECT 31.900 13.100 33.700 13.300 ;
        RECT 34.200 13.100 34.500 13.800 ;
        RECT 31.800 13.000 33.800 13.100 ;
        RECT 30.900 12.400 31.300 12.800 ;
        RECT 31.800 11.100 32.200 13.000 ;
        RECT 33.400 11.100 33.800 13.000 ;
        RECT 34.200 11.100 34.600 13.100 ;
        RECT 35.000 11.100 35.400 19.900 ;
        RECT 37.900 16.300 38.300 19.900 ;
        RECT 37.400 15.900 38.300 16.300 ;
        RECT 39.400 16.800 39.800 17.200 ;
        RECT 39.400 16.200 39.700 16.800 ;
        RECT 40.100 16.200 40.500 19.900 ;
        RECT 39.000 15.900 39.700 16.200 ;
        RECT 40.000 15.900 40.500 16.200 ;
        RECT 42.200 15.900 42.600 19.900 ;
        RECT 43.800 17.900 44.200 19.900 ;
        RECT 37.500 14.200 37.800 15.900 ;
        RECT 39.000 15.800 39.400 15.900 ;
        RECT 38.200 14.800 38.600 15.600 ;
        RECT 39.000 14.800 39.400 15.200 ;
        RECT 37.400 14.100 37.800 14.200 ;
        RECT 35.800 13.800 37.800 14.100 ;
        RECT 39.000 14.200 39.300 14.800 ;
        RECT 40.000 14.200 40.300 15.900 ;
        RECT 42.200 15.200 42.500 15.900 ;
        RECT 43.800 15.800 44.100 17.900 ;
        RECT 45.700 16.300 46.100 19.900 ;
        RECT 45.700 15.900 46.600 16.300 ;
        RECT 49.100 15.900 50.100 19.900 ;
        RECT 51.800 19.600 53.800 19.900 ;
        RECT 51.800 15.900 52.200 19.600 ;
        RECT 52.600 15.900 53.000 19.300 ;
        RECT 53.400 16.200 53.800 19.600 ;
        RECT 55.000 16.200 55.400 19.900 ;
        RECT 56.900 17.200 57.300 19.900 ;
        RECT 59.800 17.900 60.200 19.900 ;
        RECT 56.200 16.800 56.600 17.200 ;
        RECT 56.900 16.800 57.800 17.200 ;
        RECT 56.200 16.200 56.500 16.800 ;
        RECT 56.900 16.200 57.300 16.800 ;
        RECT 53.400 15.900 55.400 16.200 ;
        RECT 55.800 15.900 56.500 16.200 ;
        RECT 56.800 15.900 57.300 16.200 ;
        RECT 42.900 15.500 44.100 15.800 ;
        RECT 40.600 14.400 41.000 15.200 ;
        RECT 42.200 14.800 42.600 15.200 ;
        RECT 39.000 13.800 40.300 14.200 ;
        RECT 41.400 14.100 41.800 14.200 ;
        RECT 41.000 13.800 41.800 14.100 ;
        RECT 35.800 13.200 36.100 13.800 ;
        RECT 35.800 12.400 36.200 13.200 ;
        RECT 37.500 12.100 37.800 13.800 ;
        RECT 39.100 13.100 39.400 13.800 ;
        RECT 41.000 13.600 41.400 13.800 ;
        RECT 39.900 13.100 41.700 13.300 ;
        RECT 42.200 13.100 42.500 14.800 ;
        RECT 42.900 13.800 43.200 15.500 ;
        RECT 43.800 14.800 44.200 15.200 ;
        RECT 45.400 14.800 45.800 15.600 ;
        RECT 43.800 14.400 44.100 14.800 ;
        RECT 43.600 14.000 44.200 14.400 ;
        RECT 44.600 13.800 45.000 14.600 ;
        RECT 46.200 14.200 46.500 15.900 ;
        RECT 48.600 14.400 49.000 15.200 ;
        RECT 49.400 14.200 49.700 15.900 ;
        RECT 52.700 15.600 53.000 15.900 ;
        RECT 55.800 15.800 56.200 15.900 ;
        RECT 50.200 14.400 50.600 15.200 ;
        RECT 51.800 14.800 52.200 15.600 ;
        RECT 52.700 15.300 53.700 15.600 ;
        RECT 53.400 15.200 53.700 15.300 ;
        RECT 54.600 15.200 55.000 15.400 ;
        RECT 53.400 14.800 53.800 15.200 ;
        RECT 54.600 14.900 55.400 15.200 ;
        RECT 55.000 14.800 55.400 14.900 ;
        RECT 46.200 14.100 46.600 14.200 ;
        RECT 45.400 13.800 46.600 14.100 ;
        RECT 47.800 14.100 48.200 14.200 ;
        RECT 49.400 14.100 49.800 14.200 ;
        RECT 47.800 13.800 48.600 14.100 ;
        RECT 49.400 13.800 50.600 14.100 ;
        RECT 51.000 13.800 51.400 14.600 ;
        RECT 52.700 14.400 53.100 14.800 ;
        RECT 52.700 14.200 53.000 14.400 ;
        RECT 52.600 13.800 53.000 14.200 ;
        RECT 42.800 13.700 43.200 13.800 ;
        RECT 42.800 13.500 44.300 13.700 ;
        RECT 42.800 13.400 44.900 13.500 ;
        RECT 44.000 13.200 44.900 13.400 ;
        RECT 44.600 13.100 44.900 13.200 ;
        RECT 45.400 13.200 45.700 13.800 ;
        RECT 37.400 11.100 37.800 12.100 ;
        RECT 39.000 11.100 39.400 13.100 ;
        RECT 39.800 13.000 41.800 13.100 ;
        RECT 39.800 11.100 40.200 13.000 ;
        RECT 41.400 11.100 41.800 13.000 ;
        RECT 42.200 12.600 42.900 13.100 ;
        RECT 42.500 12.200 42.900 12.600 ;
        RECT 42.200 11.800 42.900 12.200 ;
        RECT 42.500 11.100 42.900 11.800 ;
        RECT 44.600 11.100 45.000 13.100 ;
        RECT 45.400 12.800 45.800 13.200 ;
        RECT 46.200 12.100 46.500 13.800 ;
        RECT 48.200 13.600 48.600 13.800 ;
        RECT 47.000 12.400 47.400 13.200 ;
        RECT 47.900 13.100 49.700 13.300 ;
        RECT 50.300 13.100 50.600 13.800 ;
        RECT 53.400 13.100 53.700 14.800 ;
        RECT 54.200 13.800 54.600 14.600 ;
        RECT 56.800 14.200 57.100 15.900 ;
        RECT 59.900 15.800 60.200 17.900 ;
        RECT 61.400 15.900 61.800 19.900 ;
        RECT 65.100 16.200 65.500 19.900 ;
        RECT 65.800 16.800 66.200 17.200 ;
        RECT 65.900 16.200 66.200 16.800 ;
        RECT 67.000 16.200 67.400 19.900 ;
        RECT 68.600 19.600 70.600 19.900 ;
        RECT 68.600 16.200 69.000 19.600 ;
        RECT 65.100 15.900 65.600 16.200 ;
        RECT 65.900 15.900 66.600 16.200 ;
        RECT 67.000 15.900 69.000 16.200 ;
        RECT 69.400 15.900 69.800 19.300 ;
        RECT 70.200 15.900 70.600 19.600 ;
        RECT 59.900 15.500 61.100 15.800 ;
        RECT 57.400 15.100 57.800 15.200 ;
        RECT 58.200 15.100 58.600 15.200 ;
        RECT 57.400 14.800 58.600 15.100 ;
        RECT 59.800 14.800 60.200 15.200 ;
        RECT 57.400 14.400 57.800 14.800 ;
        RECT 55.800 13.800 57.100 14.200 ;
        RECT 58.200 14.100 58.600 14.200 ;
        RECT 57.800 13.800 58.600 14.100 ;
        RECT 59.000 13.800 59.400 14.600 ;
        RECT 59.900 14.400 60.200 14.800 ;
        RECT 59.800 14.000 60.400 14.400 ;
        RECT 60.800 13.800 61.100 15.500 ;
        RECT 61.500 15.200 61.800 15.900 ;
        RECT 61.400 14.800 61.800 15.200 ;
        RECT 63.000 15.100 63.400 15.200 ;
        RECT 64.600 15.100 65.000 15.200 ;
        RECT 63.000 14.800 65.000 15.100 ;
        RECT 55.900 13.100 56.200 13.800 ;
        RECT 57.800 13.600 58.200 13.800 ;
        RECT 60.800 13.700 61.200 13.800 ;
        RECT 59.700 13.500 61.200 13.700 ;
        RECT 59.100 13.400 61.200 13.500 ;
        RECT 56.700 13.100 58.500 13.300 ;
        RECT 59.100 13.200 60.000 13.400 ;
        RECT 59.100 13.100 59.400 13.200 ;
        RECT 61.500 13.100 61.800 14.800 ;
        RECT 64.600 14.400 65.000 14.800 ;
        RECT 65.300 14.200 65.600 15.900 ;
        RECT 66.200 15.800 66.600 15.900 ;
        RECT 69.400 15.600 69.700 15.900 ;
        RECT 71.000 15.600 71.400 19.900 ;
        RECT 73.100 16.200 73.500 19.900 ;
        RECT 74.200 16.200 74.600 19.900 ;
        RECT 75.800 16.200 76.200 19.900 ;
        RECT 73.100 15.900 73.800 16.200 ;
        RECT 74.200 15.900 76.200 16.200 ;
        RECT 76.600 15.900 77.000 19.900 ;
        RECT 78.700 16.200 79.100 19.900 ;
        RECT 79.400 16.800 79.800 17.200 ;
        RECT 79.500 16.200 79.800 16.800 ;
        RECT 78.700 15.900 79.200 16.200 ;
        RECT 79.500 15.900 80.200 16.200 ;
        RECT 67.400 15.200 67.800 15.400 ;
        RECT 68.700 15.300 69.700 15.600 ;
        RECT 68.700 15.200 69.000 15.300 ;
        RECT 67.000 14.900 67.800 15.200 ;
        RECT 67.000 14.800 67.400 14.900 ;
        RECT 68.600 14.800 69.000 15.200 ;
        RECT 70.200 14.800 70.600 15.600 ;
        RECT 71.000 15.400 73.000 15.600 ;
        RECT 71.000 15.300 73.100 15.400 ;
        RECT 72.700 15.000 73.100 15.300 ;
        RECT 73.500 15.200 73.800 15.900 ;
        RECT 74.600 15.200 75.000 15.400 ;
        RECT 76.600 15.200 76.900 15.900 ;
        RECT 78.900 15.200 79.200 15.900 ;
        RECT 79.800 15.800 80.200 15.900 ;
        RECT 80.600 15.900 81.000 19.900 ;
        RECT 82.200 17.900 82.600 19.900 ;
        RECT 80.600 15.200 80.900 15.900 ;
        RECT 82.200 15.800 82.500 17.900 ;
        RECT 83.000 16.800 83.400 17.200 ;
        RECT 83.000 16.100 83.300 16.800 ;
        RECT 83.800 16.100 84.200 19.900 ;
        RECT 83.000 15.800 84.200 16.100 ;
        RECT 81.300 15.500 82.500 15.800 ;
        RECT 63.800 14.100 64.200 14.200 ;
        RECT 63.800 13.800 64.600 14.100 ;
        RECT 65.300 13.800 66.600 14.200 ;
        RECT 67.800 13.800 68.200 14.600 ;
        RECT 64.200 13.600 64.600 13.800 ;
        RECT 63.900 13.100 65.700 13.300 ;
        RECT 66.200 13.100 66.500 13.800 ;
        RECT 68.700 13.100 69.000 14.800 ;
        RECT 69.300 14.400 69.700 14.800 ;
        RECT 69.400 14.200 69.700 14.400 ;
        RECT 72.000 14.200 72.400 14.600 ;
        RECT 69.400 13.800 69.800 14.200 ;
        RECT 71.800 13.800 72.300 14.200 ;
        RECT 72.800 13.500 73.100 15.000 ;
        RECT 73.400 14.800 73.800 15.200 ;
        RECT 74.200 14.900 75.000 15.200 ;
        RECT 75.800 14.900 77.000 15.200 ;
        RECT 74.200 14.800 74.600 14.900 ;
        RECT 71.900 13.200 73.100 13.500 ;
        RECT 47.800 13.000 49.800 13.100 ;
        RECT 46.200 11.100 46.600 12.100 ;
        RECT 47.800 11.100 48.200 13.000 ;
        RECT 49.400 11.400 49.800 13.000 ;
        RECT 50.200 11.700 50.600 13.100 ;
        RECT 51.000 11.400 51.400 13.100 ;
        RECT 49.400 11.100 51.400 11.400 ;
        RECT 53.100 11.100 53.900 13.100 ;
        RECT 55.800 11.100 56.200 13.100 ;
        RECT 56.600 13.000 58.600 13.100 ;
        RECT 56.600 11.100 57.000 13.000 ;
        RECT 58.200 11.100 58.600 13.000 ;
        RECT 59.000 11.100 59.400 13.100 ;
        RECT 61.100 12.600 61.800 13.100 ;
        RECT 63.800 13.000 65.800 13.100 ;
        RECT 61.100 12.100 61.500 12.600 ;
        RECT 63.000 12.100 63.400 12.200 ;
        RECT 61.100 11.800 63.400 12.100 ;
        RECT 61.100 11.100 61.500 11.800 ;
        RECT 63.800 11.100 64.200 13.000 ;
        RECT 65.400 11.100 65.800 13.000 ;
        RECT 66.200 11.100 66.600 13.100 ;
        RECT 68.500 11.100 69.300 13.100 ;
        RECT 71.000 12.400 71.400 13.200 ;
        RECT 71.900 12.100 72.200 13.200 ;
        RECT 73.500 13.100 73.800 14.800 ;
        RECT 75.000 13.800 75.400 14.600 ;
        RECT 71.800 11.100 72.200 12.100 ;
        RECT 73.400 11.100 73.800 13.100 ;
        RECT 75.800 13.100 76.100 14.900 ;
        RECT 76.600 14.800 77.000 14.900 ;
        RECT 78.200 14.400 78.600 15.200 ;
        RECT 78.900 14.800 79.400 15.200 ;
        RECT 79.800 15.100 80.200 15.200 ;
        RECT 80.600 15.100 81.000 15.200 ;
        RECT 79.800 14.800 81.000 15.100 ;
        RECT 78.900 14.200 79.200 14.800 ;
        RECT 77.400 14.100 77.800 14.200 ;
        RECT 77.400 13.800 78.200 14.100 ;
        RECT 78.900 13.800 80.200 14.200 ;
        RECT 77.800 13.600 78.200 13.800 ;
        RECT 75.800 11.100 76.200 13.100 ;
        RECT 76.600 12.800 77.000 13.200 ;
        RECT 77.500 13.100 79.300 13.300 ;
        RECT 79.800 13.100 80.100 13.800 ;
        RECT 80.600 13.100 80.900 14.800 ;
        RECT 81.300 13.800 81.600 15.500 ;
        RECT 82.200 14.800 82.600 15.200 ;
        RECT 82.200 14.400 82.500 14.800 ;
        RECT 82.000 14.100 82.500 14.400 ;
        RECT 82.000 14.000 82.400 14.100 ;
        RECT 83.000 13.800 83.400 14.600 ;
        RECT 81.200 13.700 81.600 13.800 ;
        RECT 81.200 13.500 82.700 13.700 ;
        RECT 81.200 13.400 83.300 13.500 ;
        RECT 82.400 13.200 83.300 13.400 ;
        RECT 83.000 13.100 83.300 13.200 ;
        RECT 77.400 13.000 79.400 13.100 ;
        RECT 76.500 12.400 76.900 12.800 ;
        RECT 77.400 11.100 77.800 13.000 ;
        RECT 79.000 11.100 79.400 13.000 ;
        RECT 79.800 11.100 80.200 13.100 ;
        RECT 80.600 12.600 81.300 13.100 ;
        RECT 80.900 11.100 81.300 12.600 ;
        RECT 83.000 11.100 83.400 13.100 ;
        RECT 83.800 11.100 84.200 15.800 ;
        RECT 84.600 12.400 85.000 13.200 ;
        RECT 85.400 11.100 85.800 19.900 ;
        RECT 2.200 7.600 2.600 9.900 ;
        RECT 3.000 7.900 3.400 9.900 ;
        RECT 5.200 8.100 6.000 9.900 ;
        RECT 3.000 7.600 4.100 7.900 ;
        RECT 4.600 7.700 5.400 7.800 ;
        RECT 1.500 7.300 2.600 7.600 ;
        RECT 3.700 7.500 4.100 7.600 ;
        RECT 4.400 7.400 5.400 7.700 ;
        RECT 1.500 5.800 1.800 7.300 ;
        RECT 4.400 7.200 4.700 7.400 ;
        RECT 3.000 6.900 4.700 7.200 ;
        RECT 3.000 6.800 3.800 6.900 ;
        RECT 5.000 6.700 5.400 7.100 ;
        RECT 2.200 5.800 2.600 6.600 ;
        RECT 5.000 6.400 5.300 6.700 ;
        RECT 4.000 6.100 5.300 6.400 ;
        RECT 5.700 6.400 6.000 8.100 ;
        RECT 7.800 7.900 8.200 9.900 ;
        RECT 8.600 8.000 9.000 9.900 ;
        RECT 10.200 8.000 10.600 9.900 ;
        RECT 8.600 7.900 10.600 8.000 ;
        RECT 11.000 7.900 11.400 9.900 ;
        RECT 12.100 8.400 12.500 9.900 ;
        RECT 11.800 7.900 12.500 8.400 ;
        RECT 14.200 7.900 14.600 9.900 ;
        RECT 15.000 7.900 15.400 9.900 ;
        RECT 17.200 9.200 18.000 9.900 ;
        RECT 17.200 8.800 18.600 9.200 ;
        RECT 17.200 8.100 18.000 8.800 ;
        RECT 6.300 7.400 6.700 7.800 ;
        RECT 7.000 7.600 8.200 7.900 ;
        RECT 8.700 7.700 10.500 7.900 ;
        RECT 7.000 7.500 7.400 7.600 ;
        RECT 6.400 7.200 6.700 7.400 ;
        RECT 9.000 7.200 9.400 7.400 ;
        RECT 11.000 7.200 11.300 7.900 ;
        RECT 6.400 6.800 6.800 7.200 ;
        RECT 7.400 6.800 8.200 7.200 ;
        RECT 8.600 6.900 9.400 7.200 ;
        RECT 8.600 6.800 9.000 6.900 ;
        RECT 10.100 6.800 11.400 7.200 ;
        RECT 5.700 6.200 6.200 6.400 ;
        RECT 5.700 6.100 6.600 6.200 ;
        RECT 9.400 6.100 9.800 6.600 ;
        RECT 4.000 6.000 4.400 6.100 ;
        RECT 5.900 5.800 9.800 6.100 ;
        RECT 10.100 6.100 10.400 6.800 ;
        RECT 11.800 6.200 12.100 7.900 ;
        RECT 14.200 7.800 14.500 7.900 ;
        RECT 13.600 7.600 14.500 7.800 ;
        RECT 15.000 7.600 16.100 7.900 ;
        RECT 12.400 7.500 14.500 7.600 ;
        RECT 15.700 7.500 16.100 7.600 ;
        RECT 12.400 7.300 13.900 7.500 ;
        RECT 12.400 7.200 12.800 7.300 ;
        RECT 11.000 6.100 11.400 6.200 ;
        RECT 10.100 5.800 11.400 6.100 ;
        RECT 11.800 5.800 12.200 6.200 ;
        RECT 1.200 5.400 1.800 5.800 ;
        RECT 5.100 5.700 5.500 5.800 ;
        RECT 1.500 5.100 1.800 5.400 ;
        RECT 3.800 5.400 5.500 5.700 ;
        RECT 3.800 5.100 4.100 5.400 ;
        RECT 5.900 5.100 6.200 5.800 ;
        RECT 10.100 5.100 10.400 5.800 ;
        RECT 11.000 5.100 11.400 5.200 ;
        RECT 11.800 5.100 12.100 5.800 ;
        RECT 12.500 5.500 12.800 7.200 ;
        RECT 13.200 6.600 13.800 7.000 ;
        RECT 13.400 6.200 13.700 6.600 ;
        RECT 14.200 6.400 14.600 7.200 ;
        RECT 17.000 6.700 17.400 7.100 ;
        RECT 17.000 6.400 17.300 6.700 ;
        RECT 13.400 5.800 13.800 6.200 ;
        RECT 16.000 6.100 17.300 6.400 ;
        RECT 17.700 6.400 18.000 8.100 ;
        RECT 19.800 7.900 20.200 9.900 ;
        RECT 19.000 7.600 20.200 7.900 ;
        RECT 20.600 7.900 21.000 9.900 ;
        RECT 22.800 9.200 23.600 9.900 ;
        RECT 22.800 8.800 24.200 9.200 ;
        RECT 22.800 8.100 23.600 8.800 ;
        RECT 20.600 7.600 21.800 7.900 ;
        RECT 19.000 7.500 19.400 7.600 ;
        RECT 21.400 7.500 21.800 7.600 ;
        RECT 22.100 7.400 22.500 7.800 ;
        RECT 22.100 7.200 22.400 7.400 ;
        RECT 22.000 6.800 22.400 7.200 ;
        RECT 22.800 7.100 23.100 8.100 ;
        RECT 25.400 7.900 25.800 9.900 ;
        RECT 29.100 9.200 29.500 9.900 ;
        RECT 28.600 8.800 29.500 9.200 ;
        RECT 29.100 8.200 29.500 8.800 ;
        RECT 23.400 7.400 24.200 7.800 ;
        RECT 24.500 7.600 25.800 7.900 ;
        RECT 28.600 7.900 29.500 8.200 ;
        RECT 24.500 7.500 24.900 7.600 ;
        RECT 22.800 6.800 23.300 7.100 ;
        RECT 17.700 6.200 18.200 6.400 ;
        RECT 23.000 6.200 23.300 6.800 ;
        RECT 17.700 6.100 18.600 6.200 ;
        RECT 16.000 6.000 16.400 6.100 ;
        RECT 17.900 5.800 18.600 6.100 ;
        RECT 23.000 5.800 23.400 6.200 ;
        RECT 24.300 6.100 24.700 6.200 ;
        RECT 23.900 5.800 24.700 6.100 ;
        RECT 17.100 5.700 17.500 5.800 ;
        RECT 12.500 5.200 13.700 5.500 ;
        RECT 1.500 4.800 2.600 5.100 ;
        RECT 2.200 1.100 2.600 4.800 ;
        RECT 3.000 4.800 4.100 5.100 ;
        RECT 3.000 1.100 3.400 4.800 ;
        RECT 3.700 4.700 4.100 4.800 ;
        RECT 5.200 4.800 6.200 5.100 ;
        RECT 7.000 4.800 8.200 5.100 ;
        RECT 5.200 1.100 6.000 4.800 ;
        RECT 7.000 4.700 7.400 4.800 ;
        RECT 7.800 1.100 8.200 4.800 ;
        RECT 9.900 4.800 10.400 5.100 ;
        RECT 10.700 4.800 12.200 5.100 ;
        RECT 9.900 1.100 10.300 4.800 ;
        RECT 10.700 4.200 11.000 4.800 ;
        RECT 10.600 3.800 11.000 4.200 ;
        RECT 11.800 1.100 12.200 4.800 ;
        RECT 13.400 3.100 13.700 5.200 ;
        RECT 15.800 5.400 17.500 5.700 ;
        RECT 15.800 5.100 16.100 5.400 ;
        RECT 17.900 5.100 18.200 5.800 ;
        RECT 23.000 5.100 23.300 5.800 ;
        RECT 23.900 5.700 24.300 5.800 ;
        RECT 15.000 4.800 16.100 5.100 ;
        RECT 13.400 1.100 13.800 3.100 ;
        RECT 15.000 1.100 15.400 4.800 ;
        RECT 15.700 4.700 16.100 4.800 ;
        RECT 17.200 4.800 18.200 5.100 ;
        RECT 19.000 4.800 20.200 5.100 ;
        RECT 17.200 1.100 18.000 4.800 ;
        RECT 19.000 4.700 19.400 4.800 ;
        RECT 19.800 1.100 20.200 4.800 ;
        RECT 20.600 4.800 21.800 5.100 ;
        RECT 20.600 1.100 21.000 4.800 ;
        RECT 21.400 4.700 21.800 4.800 ;
        RECT 22.800 1.100 23.600 5.100 ;
        RECT 24.500 4.800 25.800 5.100 ;
        RECT 24.500 4.700 24.900 4.800 ;
        RECT 25.400 1.100 25.800 4.800 ;
        RECT 28.600 1.100 29.000 7.900 ;
        RECT 31.000 6.100 31.400 9.900 ;
        RECT 31.800 7.900 32.200 9.900 ;
        RECT 33.900 9.200 34.300 9.900 ;
        RECT 33.900 8.800 34.600 9.200 ;
        RECT 33.900 8.400 34.300 8.800 ;
        RECT 33.900 7.900 34.600 8.400 ;
        RECT 31.900 7.800 32.200 7.900 ;
        RECT 31.900 7.600 32.800 7.800 ;
        RECT 31.900 7.500 34.000 7.600 ;
        RECT 32.500 7.300 34.000 7.500 ;
        RECT 29.400 5.800 31.400 6.100 ;
        RECT 29.400 5.200 29.700 5.800 ;
        RECT 29.400 4.400 29.800 5.200 ;
        RECT 31.000 1.100 31.400 5.800 ;
        RECT 33.600 7.200 34.000 7.300 ;
        RECT 33.600 5.500 33.900 7.200 ;
        RECT 34.300 6.200 34.600 7.900 ;
        RECT 36.600 7.600 37.000 9.900 ;
        RECT 37.400 7.900 37.800 9.900 ;
        RECT 38.200 8.000 38.600 9.900 ;
        RECT 39.800 8.000 40.200 9.900 ;
        RECT 38.200 7.900 40.200 8.000 ;
        RECT 34.200 5.800 34.600 6.200 ;
        RECT 35.900 7.300 37.000 7.600 ;
        RECT 35.900 5.800 36.200 7.300 ;
        RECT 37.500 7.200 37.800 7.900 ;
        RECT 38.300 7.700 40.100 7.900 ;
        RECT 39.400 7.200 39.800 7.400 ;
        RECT 37.400 6.800 38.700 7.200 ;
        RECT 39.400 7.100 40.200 7.200 ;
        RECT 40.600 7.100 41.000 9.900 ;
        RECT 41.400 7.800 41.800 8.600 ;
        RECT 42.200 7.900 42.600 9.900 ;
        RECT 43.000 8.000 43.400 9.900 ;
        RECT 44.600 8.000 45.000 9.900 ;
        RECT 45.700 8.200 46.100 9.900 ;
        RECT 43.000 7.900 45.000 8.000 ;
        RECT 42.300 7.200 42.600 7.900 ;
        RECT 43.100 7.700 44.900 7.900 ;
        RECT 45.400 7.800 46.600 8.200 ;
        RECT 47.800 7.900 48.200 9.900 ;
        RECT 48.600 8.000 49.000 9.900 ;
        RECT 50.200 8.000 50.600 9.900 ;
        RECT 52.300 9.200 52.700 9.900 ;
        RECT 52.300 8.800 53.000 9.200 ;
        RECT 52.300 8.200 52.700 8.800 ;
        RECT 48.600 7.900 50.600 8.000 ;
        RECT 51.800 7.900 52.700 8.200 ;
        RECT 44.200 7.200 44.600 7.400 ;
        RECT 39.400 6.900 41.000 7.100 ;
        RECT 39.800 6.800 41.000 6.900 ;
        RECT 36.600 6.100 37.000 6.600 ;
        RECT 38.400 6.100 38.700 6.800 ;
        RECT 36.600 5.800 38.700 6.100 ;
        RECT 39.000 5.800 39.400 6.600 ;
        RECT 32.700 5.200 33.900 5.500 ;
        RECT 32.700 3.100 33.000 5.200 ;
        RECT 34.300 5.100 34.600 5.800 ;
        RECT 35.600 5.400 36.200 5.800 ;
        RECT 32.600 1.100 33.000 3.100 ;
        RECT 34.200 1.100 34.600 5.100 ;
        RECT 35.900 5.100 36.200 5.400 ;
        RECT 37.400 5.100 37.800 5.200 ;
        RECT 38.400 5.100 38.700 5.800 ;
        RECT 35.900 4.800 37.000 5.100 ;
        RECT 37.400 4.800 38.100 5.100 ;
        RECT 38.400 4.800 38.900 5.100 ;
        RECT 36.600 1.100 37.000 4.800 ;
        RECT 37.800 4.200 38.100 4.800 ;
        RECT 37.800 3.800 38.200 4.200 ;
        RECT 38.500 1.100 38.900 4.800 ;
        RECT 40.600 1.100 41.000 6.800 ;
        RECT 41.400 6.800 41.800 7.200 ;
        RECT 42.200 6.800 43.500 7.200 ;
        RECT 44.200 6.900 45.000 7.200 ;
        RECT 44.600 6.800 45.000 6.900 ;
        RECT 41.400 6.100 41.700 6.800 ;
        RECT 43.200 6.100 43.500 6.800 ;
        RECT 41.400 5.800 43.500 6.100 ;
        RECT 43.800 5.800 44.200 6.600 ;
        RECT 42.200 5.100 42.600 5.200 ;
        RECT 43.200 5.100 43.500 5.800 ;
        RECT 42.200 4.800 42.900 5.100 ;
        RECT 43.200 4.800 43.700 5.100 ;
        RECT 42.600 4.200 42.900 4.800 ;
        RECT 42.600 3.800 43.000 4.200 ;
        RECT 43.300 1.100 43.700 4.800 ;
        RECT 45.400 4.400 45.800 5.200 ;
        RECT 46.200 5.100 46.600 7.800 ;
        RECT 47.000 6.800 47.400 7.600 ;
        RECT 47.900 7.200 48.200 7.900 ;
        RECT 48.700 7.700 50.500 7.900 ;
        RECT 49.800 7.200 50.200 7.400 ;
        RECT 47.800 6.800 49.100 7.200 ;
        RECT 49.800 7.100 50.600 7.200 ;
        RECT 51.000 7.100 51.400 7.600 ;
        RECT 49.800 6.900 51.400 7.100 ;
        RECT 50.200 6.800 51.400 6.900 ;
        RECT 47.800 5.100 48.200 5.200 ;
        RECT 48.800 5.100 49.100 6.800 ;
        RECT 49.400 5.800 49.800 6.600 ;
        RECT 46.200 4.800 48.500 5.100 ;
        RECT 48.800 4.800 49.300 5.100 ;
        RECT 46.200 1.100 46.600 4.800 ;
        RECT 48.200 4.200 48.500 4.800 ;
        RECT 48.200 3.800 48.600 4.200 ;
        RECT 48.900 1.100 49.300 4.800 ;
        RECT 51.800 1.100 52.200 7.900 ;
        RECT 52.600 6.800 53.000 7.200 ;
        RECT 52.600 6.100 52.900 6.800 ;
        RECT 53.400 6.100 53.800 9.900 ;
        RECT 55.300 9.200 55.700 9.900 ;
        RECT 55.300 8.800 56.200 9.200 ;
        RECT 55.300 8.200 55.700 8.800 ;
        RECT 55.300 7.900 56.200 8.200 ;
        RECT 52.600 5.800 53.800 6.100 ;
        RECT 52.600 5.100 53.000 5.200 ;
        RECT 53.400 5.100 53.800 5.800 ;
        RECT 52.600 4.800 53.800 5.100 ;
        RECT 52.600 4.400 53.000 4.800 ;
        RECT 53.400 1.100 53.800 4.800 ;
        RECT 55.800 1.100 56.200 7.900 ;
        RECT 58.200 7.100 58.600 9.900 ;
        RECT 62.200 8.900 62.600 9.900 ;
        RECT 62.300 8.100 62.600 8.900 ;
        RECT 63.800 8.100 64.200 8.600 ;
        RECT 62.200 7.800 64.200 8.100 ;
        RECT 62.300 7.200 62.600 7.800 ;
        RECT 60.600 7.100 61.000 7.200 ;
        RECT 58.200 6.800 61.000 7.100 ;
        RECT 62.200 6.800 62.600 7.200 ;
        RECT 58.200 1.100 58.600 6.800 ;
        RECT 62.300 5.100 62.600 6.800 ;
        RECT 63.000 5.400 63.400 6.200 ;
        RECT 63.800 5.100 64.200 5.200 ;
        RECT 64.600 5.100 65.000 9.900 ;
        RECT 65.400 8.000 65.800 9.900 ;
        RECT 67.000 8.000 67.400 9.900 ;
        RECT 65.400 7.900 67.400 8.000 ;
        RECT 67.800 7.900 68.200 9.900 ;
        RECT 68.600 7.900 69.000 9.900 ;
        RECT 70.800 9.200 71.600 9.900 ;
        RECT 70.800 8.800 72.200 9.200 ;
        RECT 70.800 8.100 71.600 8.800 ;
        RECT 65.500 7.700 67.300 7.900 ;
        RECT 65.800 7.200 66.200 7.400 ;
        RECT 67.800 7.200 68.100 7.900 ;
        RECT 68.600 7.600 69.700 7.900 ;
        RECT 70.200 7.700 71.000 7.800 ;
        RECT 69.300 7.500 69.700 7.600 ;
        RECT 70.000 7.400 71.000 7.700 ;
        RECT 70.000 7.200 70.300 7.400 ;
        RECT 65.400 6.900 66.200 7.200 ;
        RECT 66.900 7.100 68.200 7.200 ;
        RECT 68.600 7.100 70.300 7.200 ;
        RECT 66.900 6.900 70.300 7.100 ;
        RECT 65.400 6.800 65.800 6.900 ;
        RECT 66.900 6.800 69.400 6.900 ;
        RECT 66.200 5.800 66.600 6.600 ;
        RECT 66.900 5.100 67.200 6.800 ;
        RECT 70.600 6.700 71.000 7.100 ;
        RECT 70.600 6.400 70.900 6.700 ;
        RECT 69.600 6.100 70.900 6.400 ;
        RECT 71.300 6.400 71.600 8.100 ;
        RECT 73.400 7.900 73.800 9.900 ;
        RECT 71.900 7.400 72.300 7.800 ;
        RECT 72.600 7.600 73.800 7.900 ;
        RECT 74.200 7.900 74.600 9.900 ;
        RECT 76.400 8.100 77.200 9.900 ;
        RECT 74.200 7.600 75.300 7.900 ;
        RECT 75.800 7.700 76.600 7.800 ;
        RECT 72.600 7.500 73.000 7.600 ;
        RECT 74.900 7.500 75.300 7.600 ;
        RECT 72.000 7.200 72.300 7.400 ;
        RECT 75.600 7.400 76.600 7.700 ;
        RECT 75.600 7.200 75.900 7.400 ;
        RECT 72.000 6.800 72.400 7.200 ;
        RECT 73.000 6.800 73.800 7.200 ;
        RECT 74.200 6.900 75.900 7.200 ;
        RECT 74.200 6.800 75.000 6.900 ;
        RECT 76.200 6.700 76.600 7.100 ;
        RECT 76.200 6.400 76.500 6.700 ;
        RECT 71.300 6.200 71.800 6.400 ;
        RECT 71.300 6.100 72.200 6.200 ;
        RECT 69.600 6.000 70.000 6.100 ;
        RECT 71.500 5.800 72.200 6.100 ;
        RECT 75.200 6.100 76.500 6.400 ;
        RECT 76.900 6.400 77.200 8.100 ;
        RECT 79.000 7.900 79.400 9.900 ;
        RECT 77.500 7.400 77.900 7.800 ;
        RECT 78.200 7.600 79.400 7.900 ;
        RECT 79.800 7.800 80.200 8.600 ;
        RECT 78.200 7.500 78.600 7.600 ;
        RECT 77.600 7.200 77.900 7.400 ;
        RECT 77.600 6.800 78.000 7.200 ;
        RECT 78.600 6.800 79.400 7.200 ;
        RECT 76.900 6.200 77.400 6.400 ;
        RECT 76.900 6.100 77.800 6.200 ;
        RECT 79.000 6.100 79.400 6.200 ;
        RECT 75.200 6.000 75.600 6.100 ;
        RECT 77.100 5.800 79.400 6.100 ;
        RECT 80.600 6.100 81.000 9.900 ;
        RECT 81.400 8.000 81.800 9.900 ;
        RECT 83.000 8.000 83.400 9.900 ;
        RECT 81.400 7.900 83.400 8.000 ;
        RECT 83.800 7.900 84.200 9.900 ;
        RECT 81.500 7.700 83.300 7.900 ;
        RECT 81.800 7.200 82.200 7.400 ;
        RECT 83.800 7.200 84.100 7.900 ;
        RECT 84.600 7.600 85.000 9.900 ;
        RECT 84.600 7.300 85.700 7.600 ;
        RECT 81.400 6.900 82.200 7.200 ;
        RECT 81.400 6.800 81.800 6.900 ;
        RECT 82.900 6.800 84.200 7.200 ;
        RECT 82.200 6.100 82.600 6.600 ;
        RECT 80.600 5.800 82.600 6.100 ;
        RECT 82.900 6.100 83.200 6.800 ;
        RECT 84.600 6.100 85.000 6.600 ;
        RECT 82.900 5.800 85.000 6.100 ;
        RECT 85.400 5.800 85.700 7.300 ;
        RECT 70.700 5.700 71.100 5.800 ;
        RECT 69.400 5.400 71.100 5.700 ;
        RECT 67.800 5.100 68.200 5.200 ;
        RECT 69.400 5.100 69.700 5.400 ;
        RECT 71.500 5.100 71.800 5.800 ;
        RECT 76.300 5.700 76.700 5.800 ;
        RECT 75.000 5.400 76.700 5.700 ;
        RECT 75.000 5.100 75.300 5.400 ;
        RECT 77.100 5.100 77.400 5.800 ;
        RECT 62.200 4.700 63.100 5.100 ;
        RECT 63.800 4.800 65.000 5.100 ;
        RECT 62.700 1.100 63.100 4.700 ;
        RECT 64.600 1.100 65.000 4.800 ;
        RECT 66.700 4.800 67.200 5.100 ;
        RECT 67.500 4.800 68.200 5.100 ;
        RECT 68.600 4.800 69.700 5.100 ;
        RECT 66.700 1.100 67.100 4.800 ;
        RECT 67.500 4.200 67.800 4.800 ;
        RECT 67.400 3.800 67.800 4.200 ;
        RECT 68.600 1.100 69.000 4.800 ;
        RECT 69.300 4.700 69.700 4.800 ;
        RECT 70.800 4.800 71.800 5.100 ;
        RECT 72.600 4.800 73.800 5.100 ;
        RECT 70.800 1.100 71.600 4.800 ;
        RECT 72.600 4.700 73.000 4.800 ;
        RECT 73.400 1.100 73.800 4.800 ;
        RECT 74.200 4.800 75.300 5.100 ;
        RECT 74.200 1.100 74.600 4.800 ;
        RECT 74.900 4.700 75.300 4.800 ;
        RECT 76.400 4.800 77.400 5.100 ;
        RECT 78.200 4.800 79.400 5.100 ;
        RECT 76.400 1.100 77.200 4.800 ;
        RECT 78.200 4.700 78.600 4.800 ;
        RECT 79.000 1.100 79.400 4.800 ;
        RECT 80.600 1.100 81.000 5.800 ;
        RECT 82.900 5.100 83.200 5.800 ;
        RECT 85.400 5.400 86.000 5.800 ;
        RECT 83.800 5.100 84.200 5.200 ;
        RECT 85.400 5.100 85.700 5.400 ;
        RECT 82.700 4.800 83.200 5.100 ;
        RECT 83.500 4.800 84.200 5.100 ;
        RECT 84.600 4.800 85.700 5.100 ;
        RECT 82.700 1.100 83.100 4.800 ;
        RECT 83.500 4.200 83.800 4.800 ;
        RECT 83.400 3.800 83.800 4.200 ;
        RECT 84.600 1.100 85.000 4.800 ;
      LAYER via1 ;
        RECT 1.400 61.800 1.800 62.200 ;
        RECT 7.000 66.800 7.400 67.200 ;
        RECT 7.800 61.800 8.200 62.200 ;
        RECT 18.200 66.800 18.600 67.200 ;
        RECT 11.000 65.800 11.400 66.200 ;
        RECT 13.400 65.800 13.800 66.200 ;
        RECT 12.600 64.800 13.000 65.200 ;
        RECT 26.200 66.800 26.600 67.200 ;
        RECT 23.800 65.800 24.200 66.200 ;
        RECT 14.200 61.800 14.600 62.200 ;
        RECT 25.400 61.800 25.800 62.200 ;
        RECT 37.400 66.800 37.800 67.200 ;
        RECT 31.800 65.800 32.200 66.200 ;
        RECT 35.000 61.800 35.400 62.200 ;
        RECT 38.200 64.800 38.600 65.200 ;
        RECT 41.400 64.800 41.800 65.200 ;
        RECT 43.000 66.800 43.400 67.200 ;
        RECT 49.400 65.800 49.800 66.200 ;
        RECT 52.600 65.800 53.000 66.200 ;
        RECT 53.400 65.800 53.800 66.200 ;
        RECT 67.000 66.800 67.400 67.200 ;
        RECT 43.000 61.800 43.400 62.200 ;
        RECT 55.800 61.800 56.200 62.200 ;
        RECT 61.400 63.800 61.800 64.200 ;
        RECT 67.800 64.800 68.200 65.200 ;
        RECT 71.000 61.800 71.400 62.200 ;
        RECT 74.200 64.800 74.600 65.200 ;
        RECT 75.000 64.800 75.400 65.200 ;
        RECT 80.600 65.800 81.000 66.200 ;
        RECT 80.600 61.800 81.000 62.200 ;
        RECT 82.200 61.800 82.600 62.200 ;
        RECT 2.200 54.800 2.600 55.200 ;
        RECT 3.000 51.800 3.400 52.200 ;
        RECT 18.200 54.800 18.600 55.200 ;
        RECT 5.400 51.800 5.800 52.200 ;
        RECT 7.800 51.800 8.200 52.200 ;
        RECT 11.000 51.800 11.400 52.200 ;
        RECT 19.000 53.800 19.400 54.200 ;
        RECT 16.600 51.800 17.000 52.200 ;
        RECT 28.700 55.900 29.100 56.300 ;
        RECT 34.200 58.800 34.600 59.200 ;
        RECT 29.300 54.900 29.700 55.300 ;
        RECT 23.000 53.800 23.400 54.200 ;
        RECT 26.200 53.800 26.600 54.200 ;
        RECT 28.700 53.100 29.100 53.500 ;
        RECT 20.600 51.800 21.000 52.200 ;
        RECT 43.800 55.800 44.200 56.200 ;
        RECT 45.400 51.800 45.800 52.200 ;
        RECT 47.000 51.800 47.400 52.200 ;
        RECT 50.200 52.800 50.600 53.200 ;
        RECT 49.400 51.800 49.800 52.200 ;
        RECT 58.200 56.800 58.600 57.200 ;
        RECT 59.000 53.800 59.400 54.200 ;
        RECT 64.600 56.800 65.000 57.200 ;
        RECT 63.000 55.800 63.400 56.200 ;
        RECT 73.400 58.800 73.800 59.200 ;
        RECT 70.200 54.800 70.600 55.200 ;
        RECT 65.400 52.800 65.800 53.200 ;
        RECT 69.400 53.800 69.800 54.200 ;
        RECT 73.400 54.800 73.800 55.200 ;
        RECT 71.000 53.800 71.400 54.200 ;
        RECT 74.200 53.800 74.600 54.200 ;
        RECT 77.400 53.800 77.800 54.200 ;
        RECT 84.600 54.800 85.000 55.200 ;
        RECT 79.000 51.800 79.400 52.200 ;
        RECT 4.600 46.800 5.000 47.200 ;
        RECT 3.800 45.800 4.200 46.200 ;
        RECT 5.400 45.800 5.800 46.200 ;
        RECT 15.000 46.800 15.400 47.200 ;
        RECT 17.400 46.800 17.800 47.200 ;
        RECT 20.600 46.800 21.000 47.200 ;
        RECT 27.800 44.800 28.200 45.200 ;
        RECT 30.200 45.800 30.600 46.200 ;
        RECT 36.600 46.800 37.000 47.200 ;
        RECT 37.400 45.800 37.800 46.200 ;
        RECT 33.400 44.800 33.800 45.200 ;
        RECT 35.000 44.800 35.400 45.200 ;
        RECT 43.000 48.800 43.400 49.200 ;
        RECT 48.600 47.800 49.000 48.200 ;
        RECT 39.000 44.800 39.400 45.200 ;
        RECT 52.600 45.800 53.000 46.200 ;
        RECT 47.800 41.800 48.200 42.200 ;
        RECT 63.800 48.800 64.200 49.200 ;
        RECT 56.600 41.800 57.000 42.200 ;
        RECT 62.200 43.800 62.600 44.200 ;
        RECT 67.800 45.800 68.200 46.200 ;
        RECT 63.800 44.800 64.200 45.200 ;
        RECT 71.000 44.800 71.400 45.200 ;
        RECT 81.400 48.800 81.800 49.200 ;
        RECT 77.400 47.800 77.800 48.200 ;
        RECT 75.000 45.800 75.400 46.200 ;
        RECT 78.200 45.800 78.600 46.200 ;
        RECT 69.400 41.800 69.800 42.200 ;
        RECT 75.000 42.800 75.400 43.200 ;
        RECT 85.400 46.800 85.800 47.200 ;
        RECT 81.400 44.800 81.800 45.200 ;
        RECT 84.600 45.800 85.000 46.200 ;
        RECT 82.200 41.800 82.600 42.200 ;
        RECT 85.400 44.800 85.800 45.200 ;
        RECT 1.300 35.900 1.700 36.300 ;
        RECT 6.200 34.800 6.600 35.200 ;
        RECT 1.300 33.100 1.700 33.500 ;
        RECT 7.800 34.800 8.200 35.200 ;
        RECT 8.600 33.800 9.000 34.200 ;
        RECT 9.400 33.800 9.800 34.200 ;
        RECT 6.200 31.800 6.600 32.200 ;
        RECT 11.000 31.800 11.400 32.200 ;
        RECT 15.000 32.800 15.400 33.200 ;
        RECT 14.200 31.800 14.600 32.200 ;
        RECT 19.800 31.800 20.200 32.200 ;
        RECT 22.200 31.800 22.600 32.200 ;
        RECT 28.600 34.800 29.000 35.200 ;
        RECT 26.200 32.800 26.600 33.200 ;
        RECT 30.200 32.800 30.600 33.200 ;
        RECT 40.600 33.800 41.000 34.200 ;
        RECT 31.800 31.800 32.200 32.200 ;
        RECT 45.400 32.800 45.800 33.200 ;
        RECT 55.800 36.800 56.200 37.200 ;
        RECT 50.200 32.800 50.600 33.200 ;
        RECT 54.200 34.800 54.600 35.200 ;
        RECT 55.800 34.800 56.200 35.200 ;
        RECT 56.600 33.800 57.000 34.200 ;
        RECT 57.400 33.800 57.800 34.200 ;
        RECT 59.800 34.800 60.200 35.200 ;
        RECT 63.000 35.800 63.400 36.200 ;
        RECT 64.600 34.800 65.000 35.200 ;
        RECT 68.600 34.800 69.000 35.200 ;
        RECT 71.000 34.800 71.400 35.200 ;
        RECT 75.800 36.800 76.200 37.200 ;
        RECT 79.800 36.800 80.200 37.200 ;
        RECT 72.600 33.800 73.000 34.200 ;
        RECT 58.200 31.800 58.600 32.200 ;
        RECT 68.600 32.800 69.000 33.200 ;
        RECT 77.400 35.800 77.800 36.200 ;
        RECT 76.600 34.800 77.000 35.200 ;
        RECT 82.200 34.800 82.600 35.200 ;
        RECT 84.600 34.800 85.000 35.200 ;
        RECT 80.600 33.800 81.000 34.200 ;
        RECT 7.000 28.800 7.400 29.200 ;
        RECT 3.800 21.800 4.200 22.200 ;
        RECT 6.200 24.800 6.600 25.200 ;
        RECT 35.000 28.800 35.400 29.200 ;
        RECT 10.200 25.800 10.600 26.200 ;
        RECT 15.000 25.800 15.400 26.200 ;
        RECT 9.400 21.800 9.800 22.200 ;
        RECT 14.200 24.800 14.600 25.200 ;
        RECT 16.600 25.800 17.000 26.200 ;
        RECT 19.800 24.800 20.200 25.200 ;
        RECT 38.200 26.800 38.600 27.200 ;
        RECT 39.000 25.800 39.400 26.200 ;
        RECT 35.000 24.800 35.400 25.200 ;
        RECT 43.000 26.800 43.400 27.200 ;
        RECT 41.400 25.800 41.800 26.200 ;
        RECT 49.400 26.800 49.800 27.200 ;
        RECT 36.600 21.800 37.000 22.200 ;
        RECT 47.800 24.800 48.200 25.200 ;
        RECT 44.600 21.800 45.000 22.200 ;
        RECT 51.800 23.800 52.200 24.200 ;
        RECT 56.600 25.800 57.000 26.200 ;
        RECT 72.600 28.800 73.000 29.200 ;
        RECT 65.400 26.800 65.800 27.200 ;
        RECT 61.400 25.800 61.800 26.200 ;
        RECT 52.600 21.800 53.000 22.200 ;
        RECT 55.800 21.800 56.200 22.200 ;
        RECT 59.000 24.800 59.400 25.200 ;
        RECT 69.400 25.800 69.800 26.200 ;
        RECT 66.200 24.800 66.600 25.200 ;
        RECT 67.000 24.800 67.400 25.200 ;
        RECT 69.400 24.800 69.800 25.200 ;
        RECT 77.400 28.800 77.800 29.200 ;
        RECT 76.600 26.800 77.000 27.200 ;
        RECT 79.000 27.800 79.400 28.200 ;
        RECT 82.200 26.800 82.600 27.200 ;
        RECT 79.800 24.800 80.200 25.200 ;
        RECT 83.000 24.800 83.400 25.200 ;
        RECT 84.600 21.800 85.000 22.200 ;
        RECT 3.800 16.800 4.200 17.200 ;
        RECT 5.400 15.800 5.800 16.200 ;
        RECT 4.600 14.800 5.000 15.200 ;
        RECT 12.600 14.800 13.000 15.200 ;
        RECT 13.400 14.800 13.800 15.200 ;
        RECT 19.000 14.800 19.400 15.200 ;
        RECT 31.000 18.800 31.400 19.200 ;
        RECT 35.000 18.800 35.400 19.200 ;
        RECT 15.000 11.800 15.400 12.200 ;
        RECT 19.800 13.800 20.200 14.200 ;
        RECT 17.400 12.800 17.800 13.200 ;
        RECT 16.600 11.800 17.000 12.200 ;
        RECT 21.400 12.800 21.800 13.200 ;
        RECT 32.600 14.800 33.000 15.200 ;
        RECT 57.400 16.800 57.800 17.200 ;
        RECT 40.600 14.800 41.000 15.200 ;
        RECT 35.800 12.800 36.200 13.200 ;
        RECT 41.400 13.800 41.800 14.200 ;
        RECT 43.800 14.000 44.200 14.400 ;
        RECT 48.600 14.800 49.000 15.200 ;
        RECT 50.200 14.800 50.600 15.200 ;
        RECT 47.000 12.800 47.400 13.200 ;
        RECT 58.200 14.800 58.600 15.200 ;
        RECT 58.200 13.800 58.600 14.200 ;
        RECT 63.000 11.800 63.400 12.200 ;
        RECT 66.200 11.800 66.600 12.200 ;
        RECT 71.000 12.800 71.400 13.200 ;
        RECT 73.400 11.800 73.800 12.200 ;
        RECT 78.200 14.800 78.600 15.200 ;
        RECT 79.000 14.800 79.400 15.200 ;
        RECT 75.800 11.800 76.200 12.200 ;
        RECT 85.400 18.800 85.800 19.200 ;
        RECT 84.600 12.800 85.000 13.200 ;
        RECT 4.600 7.400 5.000 7.800 ;
        RECT 18.200 8.800 18.600 9.200 ;
        RECT 7.800 6.800 8.200 7.200 ;
        RECT 11.000 5.800 11.400 6.200 ;
        RECT 13.400 6.600 13.800 7.000 ;
        RECT 14.200 6.800 14.600 7.200 ;
        RECT 23.800 8.800 24.200 9.200 ;
        RECT 23.800 7.400 24.200 7.800 ;
        RECT 31.000 8.800 31.400 9.200 ;
        RECT 34.200 8.800 34.600 9.200 ;
        RECT 52.600 8.800 53.000 9.200 ;
        RECT 45.400 4.800 45.800 5.200 ;
        RECT 48.600 6.800 49.000 7.200 ;
        RECT 51.000 6.800 51.400 7.200 ;
        RECT 55.800 8.800 56.200 9.200 ;
        RECT 60.600 6.800 61.000 7.200 ;
        RECT 63.000 5.800 63.400 6.200 ;
        RECT 71.800 8.800 72.200 9.200 ;
        RECT 70.200 7.400 70.600 7.800 ;
        RECT 75.800 7.400 76.200 7.800 ;
        RECT 73.400 6.800 73.800 7.200 ;
        RECT 79.000 6.800 79.400 7.200 ;
        RECT 79.000 5.800 79.400 6.200 ;
        RECT 67.800 4.800 68.200 5.200 ;
        RECT 83.800 4.800 84.200 5.200 ;
      LAYER metal2 ;
        RECT 20.600 67.800 21.000 68.200 ;
        RECT 23.800 67.800 24.200 68.200 ;
        RECT 31.800 67.800 32.200 68.200 ;
        RECT 33.400 67.800 33.800 68.200 ;
        RECT 38.200 68.100 38.600 68.200 ;
        RECT 39.000 68.100 39.400 68.200 ;
        RECT 38.200 67.800 39.400 68.100 ;
        RECT 46.200 67.800 46.600 68.200 ;
        RECT 49.400 67.800 49.800 68.200 ;
        RECT 55.000 67.800 55.400 68.200 ;
        RECT 67.000 67.800 67.400 68.200 ;
        RECT 2.200 67.100 2.600 67.200 ;
        RECT 3.000 67.100 3.400 67.200 ;
        RECT 2.200 66.800 3.400 67.100 ;
        RECT 7.000 66.800 7.400 67.200 ;
        RECT 9.400 67.100 9.800 67.200 ;
        RECT 10.200 67.100 10.600 67.200 ;
        RECT 9.400 66.800 10.600 67.100 ;
        RECT 17.400 67.100 17.800 67.200 ;
        RECT 18.200 67.100 18.600 67.200 ;
        RECT 17.400 66.800 18.600 67.100 ;
        RECT 1.400 61.800 1.800 62.200 ;
        RECT 1.400 56.200 1.700 61.800 ;
        RECT 1.400 55.800 1.800 56.200 ;
        RECT 4.600 55.800 5.000 56.200 ;
        RECT 1.400 55.100 1.800 55.200 ;
        RECT 2.200 55.100 2.600 55.200 ;
        RECT 1.400 54.800 2.600 55.100 ;
        RECT 3.000 55.100 3.400 55.200 ;
        RECT 3.800 55.100 4.200 55.200 ;
        RECT 3.000 54.800 4.200 55.100 ;
        RECT 3.000 51.800 3.400 52.200 ;
        RECT 3.000 48.200 3.300 51.800 ;
        RECT 4.600 49.200 4.900 55.800 ;
        RECT 5.400 53.800 5.800 54.200 ;
        RECT 5.400 52.200 5.700 53.800 ;
        RECT 7.000 53.200 7.300 66.800 ;
        RECT 20.600 66.200 20.900 67.800 ;
        RECT 23.800 66.200 24.100 67.800 ;
        RECT 31.800 67.200 32.100 67.800 ;
        RECT 33.400 67.200 33.700 67.800 ;
        RECT 46.200 67.200 46.500 67.800 ;
        RECT 25.400 67.100 25.800 67.200 ;
        RECT 26.200 67.100 26.600 67.200 ;
        RECT 25.400 66.800 26.600 67.100 ;
        RECT 31.800 66.800 32.200 67.200 ;
        RECT 33.400 66.800 33.800 67.200 ;
        RECT 37.400 66.800 37.800 67.200 ;
        RECT 39.000 67.100 39.400 67.200 ;
        RECT 38.200 66.800 39.400 67.100 ;
        RECT 43.000 67.100 43.400 67.200 ;
        RECT 43.800 67.100 44.200 67.200 ;
        RECT 43.000 66.800 44.200 67.100 ;
        RECT 46.200 66.800 46.600 67.200 ;
        RECT 48.600 66.800 49.000 67.200 ;
        RECT 37.400 66.200 37.700 66.800 ;
        RECT 10.200 66.100 10.600 66.200 ;
        RECT 11.000 66.100 11.400 66.200 ;
        RECT 10.200 65.800 11.400 66.100 ;
        RECT 12.600 66.100 13.000 66.200 ;
        RECT 13.400 66.100 13.800 66.200 ;
        RECT 12.600 65.800 13.800 66.100 ;
        RECT 20.600 65.800 21.000 66.200 ;
        RECT 23.800 65.800 24.200 66.200 ;
        RECT 25.400 65.800 25.800 66.200 ;
        RECT 27.000 65.800 27.400 66.200 ;
        RECT 29.400 65.800 29.800 66.200 ;
        RECT 31.000 66.100 31.400 66.200 ;
        RECT 31.800 66.100 32.200 66.200 ;
        RECT 31.000 65.800 32.200 66.100 ;
        RECT 37.400 65.800 37.800 66.200 ;
        RECT 12.600 64.800 13.000 65.200 ;
        RECT 19.000 64.800 19.400 65.200 ;
        RECT 11.000 63.800 11.400 64.200 ;
        RECT 11.000 63.200 11.300 63.800 ;
        RECT 11.000 62.800 11.400 63.200 ;
        RECT 7.800 61.800 8.200 62.200 ;
        RECT 7.800 57.200 8.100 61.800 ;
        RECT 12.600 58.200 12.900 64.800 ;
        RECT 19.000 64.200 19.300 64.800 ;
        RECT 19.000 63.800 19.400 64.200 ;
        RECT 25.400 62.200 25.700 65.800 ;
        RECT 27.000 62.200 27.300 65.800 ;
        RECT 29.400 65.200 29.700 65.800 ;
        RECT 38.200 65.200 38.500 66.800 ;
        RECT 41.400 65.800 41.800 66.200 ;
        RECT 43.800 66.100 44.200 66.200 ;
        RECT 44.600 66.100 45.000 66.200 ;
        RECT 43.800 65.800 45.000 66.100 ;
        RECT 45.400 65.800 45.800 66.200 ;
        RECT 46.200 66.100 46.600 66.200 ;
        RECT 47.000 66.100 47.400 66.200 ;
        RECT 46.200 65.800 47.400 66.100 ;
        RECT 41.400 65.200 41.700 65.800 ;
        RECT 45.400 65.200 45.700 65.800 ;
        RECT 29.400 64.800 29.800 65.200 ;
        RECT 38.200 64.800 38.600 65.200 ;
        RECT 41.400 64.800 41.800 65.200 ;
        RECT 43.800 64.800 44.200 65.200 ;
        RECT 45.400 64.800 45.800 65.200 ;
        RECT 43.800 64.200 44.100 64.800 ;
        RECT 43.800 63.800 44.200 64.200 ;
        RECT 14.200 61.800 14.600 62.200 ;
        RECT 25.400 61.800 25.800 62.200 ;
        RECT 27.000 61.800 27.400 62.200 ;
        RECT 34.200 61.800 34.600 62.200 ;
        RECT 35.000 61.800 35.400 62.200 ;
        RECT 43.000 61.800 43.400 62.200 ;
        RECT 12.600 57.800 13.000 58.200 ;
        RECT 7.800 56.800 8.200 57.200 ;
        RECT 14.200 56.200 14.500 61.800 ;
        RECT 22.200 56.800 22.600 57.200 ;
        RECT 10.200 55.800 10.600 56.200 ;
        RECT 14.200 55.800 14.600 56.200 ;
        RECT 18.200 55.800 18.600 56.200 ;
        RECT 10.200 55.200 10.500 55.800 ;
        RECT 18.200 55.200 18.500 55.800 ;
        RECT 22.200 55.200 22.500 56.800 ;
        RECT 9.400 54.800 9.800 55.200 ;
        RECT 10.200 54.800 10.600 55.200 ;
        RECT 14.200 54.800 14.600 55.200 ;
        RECT 18.200 54.800 18.600 55.200 ;
        RECT 22.200 54.800 22.600 55.200 ;
        RECT 9.400 54.200 9.700 54.800 ;
        RECT 14.200 54.200 14.500 54.800 ;
        RECT 7.800 54.100 8.200 54.200 ;
        RECT 8.600 54.100 9.000 54.200 ;
        RECT 7.800 53.800 9.000 54.100 ;
        RECT 9.400 53.800 9.800 54.200 ;
        RECT 14.200 53.800 14.600 54.200 ;
        RECT 19.000 54.100 19.400 54.200 ;
        RECT 19.800 54.100 20.200 54.200 ;
        RECT 19.000 53.800 20.200 54.100 ;
        RECT 23.000 53.800 23.400 54.200 ;
        RECT 7.000 52.800 7.400 53.200 ;
        RECT 5.400 51.800 5.800 52.200 ;
        RECT 7.800 51.800 8.200 52.200 ;
        RECT 11.000 51.800 11.400 52.200 ;
        RECT 16.600 51.800 17.000 52.200 ;
        RECT 4.600 48.800 5.000 49.200 ;
        RECT 3.000 47.800 3.400 48.200 ;
        RECT 4.600 47.200 4.900 48.800 ;
        RECT 4.600 46.800 5.000 47.200 ;
        RECT 5.400 46.200 5.700 51.800 ;
        RECT 7.800 47.100 8.100 51.800 ;
        RECT 11.000 47.200 11.300 51.800 ;
        RECT 16.600 51.200 16.900 51.800 ;
        RECT 16.600 50.800 17.000 51.200 ;
        RECT 19.000 50.200 19.300 53.800 ;
        RECT 19.800 52.800 20.200 53.200 ;
        RECT 19.800 50.200 20.100 52.800 ;
        RECT 20.600 51.800 21.000 52.200 ;
        RECT 11.800 49.800 12.200 50.200 ;
        RECT 19.000 49.800 19.400 50.200 ;
        RECT 19.800 49.800 20.200 50.200 ;
        RECT 11.800 47.200 12.100 49.800 ;
        RECT 12.600 48.800 13.000 49.200 ;
        RECT 16.600 48.800 17.000 49.200 ;
        RECT 12.600 48.200 12.900 48.800 ;
        RECT 12.600 47.800 13.000 48.200 ;
        RECT 14.200 47.800 14.600 48.200 ;
        RECT 8.600 47.100 9.000 47.200 ;
        RECT 7.800 46.800 9.000 47.100 ;
        RECT 11.000 46.800 11.400 47.200 ;
        RECT 11.800 46.800 12.200 47.200 ;
        RECT 2.200 46.100 2.600 46.200 ;
        RECT 3.000 46.100 3.400 46.200 ;
        RECT 2.200 45.800 3.400 46.100 ;
        RECT 3.800 45.800 4.200 46.200 ;
        RECT 5.400 45.800 5.800 46.200 ;
        RECT 6.200 46.100 6.600 46.200 ;
        RECT 7.000 46.100 7.400 46.200 ;
        RECT 6.200 45.800 7.400 46.100 ;
        RECT 3.800 37.200 4.100 45.800 ;
        RECT 6.200 45.100 6.600 45.200 ;
        RECT 7.000 45.100 7.400 45.200 ;
        RECT 6.200 44.800 7.400 45.100 ;
        RECT 3.800 36.800 4.200 37.200 ;
        RECT 1.300 35.900 1.700 36.300 ;
        RECT 4.600 35.900 5.000 36.300 ;
        RECT 1.300 33.500 1.600 35.900 ;
        RECT 2.600 34.200 3.000 34.300 ;
        RECT 4.700 34.200 5.000 35.900 ;
        RECT 6.200 36.100 6.600 36.200 ;
        RECT 7.000 36.100 7.400 36.200 ;
        RECT 6.200 35.800 7.400 36.100 ;
        RECT 7.800 35.800 8.200 36.200 ;
        RECT 7.800 35.200 8.100 35.800 ;
        RECT 2.600 33.900 5.000 34.200 ;
        RECT 4.700 33.500 5.000 33.900 ;
        RECT 6.200 34.800 6.600 35.200 ;
        RECT 7.800 34.800 8.200 35.200 ;
        RECT 6.200 34.200 6.500 34.800 ;
        RECT 8.600 34.200 8.900 46.800 ;
        RECT 14.200 46.200 14.500 47.800 ;
        RECT 15.000 46.800 15.400 47.200 ;
        RECT 15.800 46.800 16.200 47.200 ;
        RECT 15.000 46.200 15.300 46.800 ;
        RECT 15.800 46.200 16.100 46.800 ;
        RECT 16.600 46.200 16.900 48.800 ;
        RECT 17.400 47.800 17.800 48.200 ;
        RECT 18.200 47.800 18.600 48.200 ;
        RECT 19.000 47.800 19.400 48.200 ;
        RECT 17.400 47.200 17.700 47.800 ;
        RECT 17.400 46.800 17.800 47.200 ;
        RECT 10.200 46.100 10.600 46.200 ;
        RECT 11.000 46.100 11.400 46.200 ;
        RECT 10.200 45.800 11.400 46.100 ;
        RECT 11.800 45.800 12.200 46.200 ;
        RECT 14.200 45.800 14.600 46.200 ;
        RECT 15.000 45.800 15.400 46.200 ;
        RECT 15.800 45.800 16.200 46.200 ;
        RECT 16.600 45.800 17.000 46.200 ;
        RECT 11.800 45.200 12.100 45.800 ;
        RECT 9.400 44.800 9.800 45.200 ;
        RECT 11.800 44.800 12.200 45.200 ;
        RECT 9.400 43.200 9.700 44.800 ;
        RECT 9.400 42.800 9.800 43.200 ;
        RECT 10.200 42.800 10.600 43.200 ;
        RECT 9.400 34.800 9.800 35.200 ;
        RECT 9.400 34.200 9.700 34.800 ;
        RECT 6.200 33.800 6.600 34.200 ;
        RECT 8.600 33.800 9.000 34.200 ;
        RECT 9.400 33.800 9.800 34.200 ;
        RECT 1.300 33.100 1.700 33.500 ;
        RECT 4.600 33.100 5.000 33.500 ;
        RECT 8.600 33.200 8.900 33.800 ;
        RECT 8.600 32.800 9.000 33.200 ;
        RECT 6.200 31.800 6.600 32.200 ;
        RECT 6.200 31.200 6.500 31.800 ;
        RECT 6.200 30.800 6.600 31.200 ;
        RECT 8.600 30.800 9.000 31.200 ;
        RECT 6.200 29.100 6.600 29.200 ;
        RECT 7.000 29.100 7.400 29.200 ;
        RECT 6.200 28.800 7.400 29.100 ;
        RECT 1.500 27.800 1.900 27.900 ;
        RECT 1.500 27.500 4.300 27.800 ;
        RECT 4.600 27.500 5.000 27.900 ;
        RECT 1.500 25.100 1.800 27.500 ;
        RECT 2.200 27.400 2.600 27.500 ;
        RECT 3.900 27.400 4.300 27.500 ;
        RECT 4.700 27.100 5.000 27.500 ;
        RECT 2.200 26.800 5.000 27.100 ;
        RECT 2.200 26.100 2.500 26.800 ;
        RECT 2.100 25.700 2.500 26.100 ;
        RECT 4.700 25.100 5.000 26.800 ;
        RECT 7.800 27.800 8.200 28.200 ;
        RECT 7.800 27.200 8.100 27.800 ;
        RECT 7.800 26.800 8.200 27.200 ;
        RECT 1.500 24.700 1.900 25.100 ;
        RECT 4.600 24.700 5.000 25.100 ;
        RECT 6.200 25.100 6.600 25.200 ;
        RECT 7.000 25.100 7.400 25.200 ;
        RECT 6.200 24.800 7.400 25.100 ;
        RECT 3.800 21.800 4.200 22.200 ;
        RECT 3.800 18.200 4.100 21.800 ;
        RECT 5.400 18.800 5.800 19.200 ;
        RECT 3.800 17.800 4.200 18.200 ;
        RECT 3.800 16.800 4.200 17.200 ;
        RECT 3.800 16.200 4.100 16.800 ;
        RECT 5.400 16.200 5.700 18.800 ;
        RECT 6.200 17.800 6.600 18.200 ;
        RECT 3.800 15.800 4.200 16.200 ;
        RECT 5.400 15.800 5.800 16.200 ;
        RECT 6.200 15.200 6.500 17.800 ;
        RECT 7.000 15.800 7.400 16.200 ;
        RECT 7.000 15.200 7.300 15.800 ;
        RECT 4.600 15.100 5.000 15.200 ;
        RECT 5.400 15.100 5.800 15.200 ;
        RECT 4.600 14.800 5.800 15.100 ;
        RECT 6.200 14.800 6.600 15.200 ;
        RECT 7.000 14.800 7.400 15.200 ;
        RECT 6.200 14.100 6.600 14.200 ;
        RECT 7.000 14.100 7.400 14.200 ;
        RECT 6.200 13.800 7.400 14.100 ;
        RECT 7.800 9.200 8.100 26.800 ;
        RECT 8.600 25.200 8.900 30.800 ;
        RECT 9.400 25.200 9.700 33.800 ;
        RECT 10.200 26.200 10.500 42.800 ;
        RECT 11.800 36.200 12.100 44.800 ;
        RECT 18.200 38.200 18.500 47.800 ;
        RECT 18.200 37.800 18.600 38.200 ;
        RECT 12.600 36.800 13.000 37.200 ;
        RECT 11.000 35.800 11.400 36.200 ;
        RECT 11.800 35.800 12.200 36.200 ;
        RECT 11.000 34.200 11.300 35.800 ;
        RECT 11.800 35.200 12.100 35.800 ;
        RECT 11.800 34.800 12.200 35.200 ;
        RECT 11.000 33.800 11.400 34.200 ;
        RECT 11.800 33.800 12.200 34.200 ;
        RECT 11.800 33.200 12.100 33.800 ;
        RECT 11.800 32.800 12.200 33.200 ;
        RECT 11.000 31.800 11.400 32.200 ;
        RECT 10.200 25.800 10.600 26.200 ;
        RECT 8.600 24.800 9.000 25.200 ;
        RECT 9.400 24.800 9.800 25.200 ;
        RECT 10.200 24.100 10.600 24.200 ;
        RECT 11.000 24.100 11.300 31.800 ;
        RECT 11.800 28.800 12.200 29.200 ;
        RECT 11.800 27.200 12.100 28.800 ;
        RECT 11.800 26.800 12.200 27.200 ;
        RECT 10.200 23.800 11.300 24.100 ;
        RECT 12.600 26.200 12.900 36.800 ;
        RECT 15.800 35.100 16.200 35.200 ;
        RECT 16.600 35.100 17.000 35.200 ;
        RECT 15.800 34.800 17.000 35.100 ;
        RECT 17.400 34.100 17.800 34.200 ;
        RECT 18.200 34.100 18.500 37.800 ;
        RECT 17.400 33.800 18.500 34.100 ;
        RECT 19.000 34.200 19.300 47.800 ;
        RECT 19.800 45.200 20.100 49.800 ;
        RECT 20.600 48.200 20.900 51.800 ;
        RECT 23.000 48.200 23.300 53.800 ;
        RECT 25.400 53.200 25.700 61.800 ;
        RECT 34.200 59.200 34.500 61.800 ;
        RECT 35.000 59.200 35.300 61.800 ;
        RECT 34.200 58.800 34.600 59.200 ;
        RECT 35.000 58.800 35.400 59.200 ;
        RECT 42.200 57.800 42.600 58.200 ;
        RECT 35.800 56.800 36.200 57.200 ;
        RECT 27.000 55.800 27.400 56.200 ;
        RECT 28.700 55.900 29.100 56.300 ;
        RECT 31.800 55.900 32.200 56.300 ;
        RECT 26.200 53.800 26.600 54.200 ;
        RECT 25.400 52.800 25.800 53.200 ;
        RECT 20.600 47.800 21.000 48.200 ;
        RECT 23.000 47.800 23.400 48.200 ;
        RECT 23.000 47.200 23.300 47.800 ;
        RECT 20.600 46.800 21.000 47.200 ;
        RECT 21.400 47.100 21.800 47.200 ;
        RECT 22.200 47.100 22.600 47.200 ;
        RECT 21.400 46.800 22.600 47.100 ;
        RECT 23.000 46.800 23.400 47.200 ;
        RECT 25.400 46.800 25.800 47.200 ;
        RECT 20.600 46.200 20.900 46.800 ;
        RECT 20.600 45.800 21.000 46.200 ;
        RECT 19.800 44.800 20.200 45.200 ;
        RECT 25.400 39.200 25.700 46.800 ;
        RECT 26.200 45.200 26.500 53.800 ;
        RECT 27.000 53.200 27.300 55.800 ;
        RECT 28.700 53.500 29.000 55.900 ;
        RECT 29.300 54.900 29.700 55.300 ;
        RECT 29.400 54.200 29.700 54.900 ;
        RECT 31.900 54.200 32.200 55.900 ;
        RECT 35.800 54.200 36.100 56.800 ;
        RECT 36.600 54.800 37.000 55.200 ;
        RECT 39.000 54.800 39.400 55.200 ;
        RECT 29.400 53.900 32.200 54.200 ;
        RECT 29.400 53.500 29.800 53.600 ;
        RECT 31.100 53.500 31.500 53.600 ;
        RECT 31.900 53.500 32.200 53.900 ;
        RECT 28.700 53.200 31.500 53.500 ;
        RECT 27.000 52.800 27.400 53.200 ;
        RECT 28.700 53.100 29.100 53.200 ;
        RECT 31.800 53.100 32.200 53.500 ;
        RECT 34.200 53.800 34.600 54.200 ;
        RECT 35.800 53.800 36.200 54.200 ;
        RECT 26.200 44.800 26.600 45.200 ;
        RECT 25.400 38.800 25.800 39.200 ;
        RECT 27.000 37.200 27.300 52.800 ;
        RECT 29.400 51.800 29.800 52.200 ;
        RECT 29.400 48.200 29.700 51.800 ;
        RECT 34.200 49.200 34.500 53.800 ;
        RECT 36.600 51.200 36.900 54.800 ;
        RECT 39.000 54.200 39.300 54.800 ;
        RECT 39.000 53.800 39.400 54.200 ;
        RECT 42.200 53.100 42.500 57.800 ;
        RECT 43.000 56.200 43.300 61.800 ;
        RECT 43.800 58.800 44.200 59.200 ;
        RECT 45.400 58.800 45.800 59.200 ;
        RECT 43.800 56.200 44.100 58.800 ;
        RECT 45.400 56.200 45.700 58.800 ;
        RECT 43.000 55.800 43.400 56.200 ;
        RECT 43.800 55.800 44.200 56.200 ;
        RECT 45.400 55.800 45.800 56.200 ;
        RECT 47.000 55.100 47.400 55.200 ;
        RECT 47.800 55.100 48.200 55.200 ;
        RECT 47.000 54.800 48.200 55.100 ;
        RECT 42.200 52.800 43.300 53.100 ;
        RECT 42.200 51.800 42.600 52.200 ;
        RECT 36.600 50.800 37.000 51.200 ;
        RECT 37.400 50.800 37.800 51.200 ;
        RECT 36.600 49.800 37.000 50.200 ;
        RECT 34.200 48.800 34.600 49.200 ;
        RECT 29.400 47.800 29.800 48.200 ;
        RECT 36.600 47.200 36.900 49.800 ;
        RECT 28.600 46.800 29.000 47.200 ;
        RECT 30.200 47.100 30.600 47.200 ;
        RECT 31.000 47.100 31.400 47.200 ;
        RECT 30.200 46.800 31.400 47.100 ;
        RECT 35.000 47.100 35.400 47.200 ;
        RECT 35.800 47.100 36.200 47.200 ;
        RECT 35.000 46.800 36.200 47.100 ;
        RECT 36.600 46.800 37.000 47.200 ;
        RECT 28.600 46.200 28.900 46.800 ;
        RECT 37.400 46.200 37.700 50.800 ;
        RECT 39.800 48.800 40.200 49.200 ;
        RECT 39.800 47.200 40.100 48.800 ;
        RECT 42.200 47.200 42.500 51.800 ;
        RECT 43.000 49.200 43.300 52.800 ;
        RECT 45.400 51.800 45.800 52.200 ;
        RECT 47.000 51.800 47.400 52.200 ;
        RECT 43.000 48.800 43.400 49.200 ;
        RECT 45.400 47.200 45.700 51.800 ;
        RECT 47.000 51.200 47.300 51.800 ;
        RECT 47.000 50.800 47.400 51.200 ;
        RECT 48.600 48.200 48.900 66.800 ;
        RECT 49.400 66.200 49.700 67.800 ;
        RECT 50.200 66.800 50.600 67.200 ;
        RECT 53.400 66.800 53.800 67.200 ;
        RECT 50.200 66.200 50.500 66.800 ;
        RECT 53.400 66.200 53.700 66.800 ;
        RECT 55.000 66.200 55.300 67.800 ;
        RECT 67.000 67.200 67.300 67.800 ;
        RECT 69.300 67.500 69.700 67.900 ;
        RECT 72.600 67.500 73.000 67.900 ;
        RECT 67.000 66.800 67.400 67.200 ;
        RECT 49.400 65.800 49.800 66.200 ;
        RECT 50.200 65.800 50.600 66.200 ;
        RECT 52.600 65.800 53.000 66.200 ;
        RECT 53.400 65.800 53.800 66.200 ;
        RECT 55.000 65.800 55.400 66.200 ;
        RECT 52.600 65.200 52.900 65.800 ;
        RECT 52.600 64.800 53.000 65.200 ;
        RECT 67.800 65.100 68.200 65.200 ;
        RECT 68.600 65.100 69.000 65.200 ;
        RECT 67.800 64.800 69.000 65.100 ;
        RECT 69.300 65.100 69.600 67.500 ;
        RECT 72.700 67.100 73.000 67.500 ;
        RECT 70.600 66.800 73.000 67.100 ;
        RECT 70.600 66.700 71.000 66.800 ;
        RECT 72.700 65.100 73.000 66.800 ;
        RECT 75.800 66.800 76.200 67.200 ;
        RECT 75.000 65.800 75.400 66.200 ;
        RECT 75.000 65.200 75.300 65.800 ;
        RECT 69.300 64.700 69.700 65.100 ;
        RECT 72.600 64.700 73.000 65.100 ;
        RECT 74.200 64.800 74.600 65.200 ;
        RECT 75.000 64.800 75.400 65.200 ;
        RECT 61.400 63.800 61.800 64.200 ;
        RECT 55.800 61.800 56.200 62.200 ;
        RECT 59.800 61.800 60.200 62.200 ;
        RECT 55.800 60.200 56.100 61.800 ;
        RECT 55.800 59.800 56.200 60.200 ;
        RECT 52.600 56.800 53.000 57.200 ;
        RECT 58.200 57.100 58.600 57.200 ;
        RECT 59.000 57.100 59.400 57.200 ;
        RECT 58.200 56.800 59.400 57.100 ;
        RECT 52.600 56.200 52.900 56.800 ;
        RECT 59.800 56.200 60.100 61.800 ;
        RECT 60.600 56.800 61.000 57.200 ;
        RECT 60.600 56.200 60.900 56.800 ;
        RECT 50.200 55.800 50.600 56.200 ;
        RECT 52.600 55.800 53.000 56.200 ;
        RECT 53.400 56.100 53.800 56.200 ;
        RECT 54.200 56.100 54.600 56.200 ;
        RECT 53.400 55.800 54.600 56.100 ;
        RECT 59.800 55.800 60.200 56.200 ;
        RECT 60.600 55.800 61.000 56.200 ;
        RECT 50.200 53.200 50.500 55.800 ;
        RECT 52.600 55.100 53.000 55.200 ;
        RECT 53.400 55.100 53.800 55.200 ;
        RECT 52.600 54.800 53.800 55.100 ;
        RECT 59.000 54.800 59.400 55.200 ;
        RECT 59.800 54.800 60.200 55.200 ;
        RECT 59.000 54.200 59.300 54.800 ;
        RECT 57.400 53.800 57.800 54.200 ;
        RECT 59.000 53.800 59.400 54.200 ;
        RECT 50.200 52.800 50.600 53.200 ;
        RECT 49.400 51.800 49.800 52.200 ;
        RECT 49.400 49.200 49.700 51.800 ;
        RECT 49.400 48.800 49.800 49.200 ;
        RECT 50.200 48.200 50.500 52.800 ;
        RECT 53.400 51.800 53.800 52.200 ;
        RECT 48.600 47.800 49.000 48.200 ;
        RECT 50.200 47.800 50.600 48.200 ;
        RECT 51.800 48.100 52.200 48.200 ;
        RECT 52.600 48.100 53.000 48.200 ;
        RECT 51.800 47.800 53.000 48.100 ;
        RECT 39.800 46.800 40.200 47.200 ;
        RECT 42.200 46.800 42.600 47.200 ;
        RECT 45.400 46.800 45.800 47.200 ;
        RECT 52.600 46.800 53.000 47.200 ;
        RECT 42.200 46.200 42.500 46.800 ;
        RECT 45.400 46.200 45.700 46.800 ;
        RECT 52.600 46.200 52.900 46.800 ;
        RECT 27.800 45.800 28.200 46.200 ;
        RECT 28.600 45.800 29.000 46.200 ;
        RECT 30.200 45.800 30.600 46.200 ;
        RECT 31.000 45.800 31.400 46.200 ;
        RECT 31.800 45.800 32.200 46.200 ;
        RECT 37.400 45.800 37.800 46.200 ;
        RECT 39.000 45.800 39.400 46.200 ;
        RECT 42.200 45.800 42.600 46.200 ;
        RECT 45.400 45.800 45.800 46.200 ;
        RECT 47.000 46.100 47.400 46.200 ;
        RECT 47.800 46.100 48.200 46.200 ;
        RECT 47.000 45.800 48.200 46.100 ;
        RECT 49.400 46.100 49.800 46.200 ;
        RECT 50.200 46.100 50.600 46.200 ;
        RECT 49.400 45.800 50.600 46.100 ;
        RECT 52.600 45.800 53.000 46.200 ;
        RECT 27.800 45.200 28.100 45.800 ;
        RECT 30.200 45.200 30.500 45.800 ;
        RECT 31.000 45.200 31.300 45.800 ;
        RECT 31.800 45.200 32.100 45.800 ;
        RECT 27.800 44.800 28.200 45.200 ;
        RECT 30.200 44.800 30.600 45.200 ;
        RECT 31.000 44.800 31.400 45.200 ;
        RECT 31.800 44.800 32.200 45.200 ;
        RECT 33.400 45.100 33.800 45.200 ;
        RECT 35.000 45.100 35.400 45.200 ;
        RECT 33.400 44.800 35.400 45.100 ;
        RECT 30.200 41.800 30.600 42.200 ;
        RECT 25.400 36.800 25.800 37.200 ;
        RECT 27.000 36.800 27.400 37.200 ;
        RECT 19.800 36.100 20.200 36.200 ;
        RECT 20.600 36.100 21.000 36.200 ;
        RECT 19.800 35.800 21.000 36.100 ;
        RECT 23.800 36.100 24.200 36.200 ;
        RECT 24.600 36.100 25.000 36.200 ;
        RECT 23.800 35.800 25.000 36.100 ;
        RECT 20.600 35.200 20.900 35.800 ;
        RECT 20.600 34.800 21.000 35.200 ;
        RECT 21.400 34.800 21.800 35.200 ;
        RECT 19.000 33.800 19.400 34.200 ;
        RECT 20.600 33.800 21.000 34.200 ;
        RECT 14.200 32.800 14.600 33.200 ;
        RECT 15.000 32.800 15.400 33.200 ;
        RECT 14.200 32.200 14.500 32.800 ;
        RECT 14.200 31.800 14.600 32.200 ;
        RECT 15.000 28.200 15.300 32.800 ;
        RECT 18.200 28.800 18.600 29.200 ;
        RECT 14.200 28.100 14.600 28.200 ;
        RECT 15.000 28.100 15.400 28.200 ;
        RECT 14.200 27.800 15.400 28.100 ;
        RECT 16.600 27.800 17.000 28.200 ;
        RECT 16.600 26.200 16.900 27.800 ;
        RECT 18.200 26.200 18.500 28.800 ;
        RECT 12.600 25.800 13.000 26.200 ;
        RECT 15.000 25.800 15.400 26.200 ;
        RECT 16.600 25.800 17.000 26.200 ;
        RECT 18.200 25.800 18.600 26.200 ;
        RECT 9.400 21.800 9.800 22.200 ;
        RECT 9.400 19.200 9.700 21.800 ;
        RECT 9.400 18.800 9.800 19.200 ;
        RECT 11.000 17.800 11.400 18.200 ;
        RECT 9.400 16.800 9.800 17.200 ;
        RECT 9.400 13.200 9.700 16.800 ;
        RECT 11.000 14.200 11.300 17.800 ;
        RECT 12.600 15.200 12.900 25.800 ;
        RECT 15.000 25.200 15.300 25.800 ;
        RECT 14.200 24.800 14.600 25.200 ;
        RECT 15.000 24.800 15.400 25.200 ;
        RECT 13.400 23.800 13.800 24.200 ;
        RECT 13.400 18.200 13.700 23.800 ;
        RECT 14.200 23.200 14.500 24.800 ;
        RECT 14.200 22.800 14.600 23.200 ;
        RECT 15.000 21.800 15.400 22.200 ;
        RECT 18.200 21.800 18.600 22.200 ;
        RECT 14.200 18.800 14.600 19.200 ;
        RECT 13.400 17.800 13.800 18.200 ;
        RECT 13.400 15.200 13.700 17.800 ;
        RECT 12.600 14.800 13.000 15.200 ;
        RECT 13.400 14.800 13.800 15.200 ;
        RECT 12.600 14.200 12.900 14.800 ;
        RECT 11.000 13.800 11.400 14.200 ;
        RECT 12.600 13.800 13.000 14.200 ;
        RECT 9.400 12.800 9.800 13.200 ;
        RECT 7.800 8.800 8.200 9.200 ;
        RECT 3.000 7.800 3.400 8.200 ;
        RECT 3.000 7.200 3.300 7.800 ;
        RECT 3.700 7.500 4.100 7.900 ;
        RECT 4.600 7.500 6.700 7.800 ;
        RECT 7.000 7.500 7.400 7.900 ;
        RECT 3.000 6.800 3.400 7.200 ;
        RECT 2.200 6.100 2.600 6.200 ;
        RECT 3.000 6.100 3.400 6.200 ;
        RECT 2.200 5.800 3.400 6.100 ;
        RECT 3.700 5.100 4.000 7.500 ;
        RECT 4.600 7.400 5.000 7.500 ;
        RECT 6.300 7.400 6.700 7.500 ;
        RECT 7.100 7.100 7.400 7.500 ;
        RECT 5.000 6.800 7.400 7.100 ;
        RECT 7.800 7.200 8.100 8.800 ;
        RECT 7.800 6.800 8.200 7.200 ;
        RECT 8.600 7.100 9.000 7.200 ;
        RECT 9.400 7.100 9.700 12.800 ;
        RECT 8.600 6.800 9.700 7.100 ;
        RECT 13.400 9.800 13.800 10.200 ;
        RECT 13.400 7.000 13.700 9.800 ;
        RECT 14.200 7.200 14.500 18.800 ;
        RECT 15.000 16.200 15.300 21.800 ;
        RECT 18.200 19.200 18.500 21.800 ;
        RECT 18.200 18.800 18.600 19.200 ;
        RECT 18.200 17.800 18.600 18.200 ;
        RECT 15.000 15.800 15.400 16.200 ;
        RECT 15.800 15.100 16.200 15.200 ;
        RECT 16.600 15.100 17.000 15.200 ;
        RECT 15.800 14.800 17.000 15.100 ;
        RECT 18.200 14.200 18.500 17.800 ;
        RECT 19.000 17.200 19.300 33.800 ;
        RECT 19.800 31.800 20.200 32.200 ;
        RECT 19.800 28.200 20.100 31.800 ;
        RECT 20.600 31.200 20.900 33.800 ;
        RECT 20.600 30.800 21.000 31.200 ;
        RECT 19.800 27.800 20.200 28.200 ;
        RECT 20.600 27.800 21.000 28.200 ;
        RECT 20.600 27.200 20.900 27.800 ;
        RECT 20.600 26.800 21.000 27.200 ;
        RECT 19.800 25.800 20.200 26.200 ;
        RECT 19.800 25.200 20.100 25.800 ;
        RECT 19.800 24.800 20.200 25.200 ;
        RECT 20.600 18.200 20.900 26.800 ;
        RECT 21.400 26.200 21.700 34.800 ;
        RECT 23.000 32.800 23.400 33.200 ;
        RECT 22.200 31.800 22.600 32.200 ;
        RECT 22.200 29.200 22.500 31.800 ;
        RECT 22.200 28.800 22.600 29.200 ;
        RECT 23.000 26.200 23.300 32.800 ;
        RECT 21.400 25.800 21.800 26.200 ;
        RECT 23.000 25.800 23.400 26.200 ;
        RECT 25.400 25.200 25.700 36.800 ;
        RECT 28.600 35.800 29.000 36.200 ;
        RECT 28.600 35.200 28.900 35.800 ;
        RECT 28.600 34.800 29.000 35.200 ;
        RECT 28.600 33.800 29.000 34.200 ;
        RECT 28.600 33.200 28.900 33.800 ;
        RECT 30.200 33.200 30.500 41.800 ;
        RECT 31.000 35.800 31.400 36.200 ;
        RECT 31.000 35.200 31.300 35.800 ;
        RECT 31.000 34.800 31.400 35.200 ;
        RECT 36.600 35.100 37.000 35.200 ;
        RECT 37.400 35.100 37.700 45.800 ;
        RECT 39.000 45.200 39.300 45.800 ;
        RECT 39.000 44.800 39.400 45.200 ;
        RECT 41.400 43.100 41.800 43.200 ;
        RECT 42.200 43.100 42.600 43.200 ;
        RECT 41.400 42.800 42.600 43.100 ;
        RECT 47.800 41.800 48.200 42.200 ;
        RECT 47.800 40.200 48.100 41.800 ;
        RECT 47.800 39.800 48.200 40.200 ;
        RECT 43.000 37.800 43.400 38.200 ;
        RECT 36.600 34.800 37.700 35.100 ;
        RECT 40.600 35.800 41.000 36.200 ;
        RECT 42.200 35.800 42.600 36.200 ;
        RECT 40.600 35.200 40.900 35.800 ;
        RECT 40.600 34.800 41.000 35.200 ;
        RECT 34.200 33.800 34.600 34.200 ;
        RECT 35.800 33.800 36.200 34.200 ;
        RECT 34.200 33.200 34.500 33.800 ;
        RECT 26.200 32.800 26.600 33.200 ;
        RECT 28.600 32.800 29.000 33.200 ;
        RECT 30.200 32.800 30.600 33.200 ;
        RECT 34.200 32.800 34.600 33.200 ;
        RECT 26.200 32.200 26.500 32.800 ;
        RECT 26.200 31.800 26.600 32.200 ;
        RECT 30.200 28.200 30.500 32.800 ;
        RECT 35.800 32.200 36.100 33.800 ;
        RECT 36.600 32.800 37.000 33.200 ;
        RECT 31.800 31.800 32.200 32.200 ;
        RECT 34.200 31.800 34.600 32.200 ;
        RECT 35.800 31.800 36.200 32.200 ;
        RECT 31.800 29.200 32.100 31.800 ;
        RECT 31.800 28.800 32.200 29.200 ;
        RECT 33.400 28.800 33.800 29.200 ;
        RECT 30.200 27.800 30.600 28.200 ;
        RECT 32.600 26.800 33.000 27.200 ;
        RECT 32.600 26.200 32.900 26.800 ;
        RECT 33.400 26.200 33.700 28.800 ;
        RECT 32.600 25.800 33.000 26.200 ;
        RECT 33.400 25.800 33.800 26.200 ;
        RECT 25.400 24.800 25.800 25.200 ;
        RECT 21.400 21.800 21.800 22.200 ;
        RECT 20.600 17.800 21.000 18.200 ;
        RECT 19.000 16.800 19.400 17.200 ;
        RECT 20.600 15.800 21.000 16.200 ;
        RECT 20.600 15.200 20.900 15.800 ;
        RECT 19.000 14.800 19.400 15.200 ;
        RECT 20.600 14.800 21.000 15.200 ;
        RECT 18.200 13.800 18.600 14.200 ;
        RECT 17.400 13.100 17.800 13.200 ;
        RECT 18.200 13.100 18.600 13.200 ;
        RECT 17.400 12.800 18.600 13.100 ;
        RECT 15.000 11.800 15.400 12.200 ;
        RECT 16.600 11.800 17.000 12.200 ;
        RECT 19.000 12.100 19.300 14.800 ;
        RECT 19.800 13.800 20.200 14.200 ;
        RECT 19.800 13.200 20.100 13.800 ;
        RECT 21.400 13.200 21.700 21.800 ;
        RECT 25.400 18.200 25.700 24.800 ;
        RECT 31.000 22.800 31.400 23.200 ;
        RECT 29.400 21.800 29.800 22.200 ;
        RECT 25.400 17.800 25.800 18.200 ;
        RECT 22.200 16.800 22.600 17.200 ;
        RECT 22.200 16.200 22.500 16.800 ;
        RECT 25.400 16.200 25.700 17.800 ;
        RECT 22.200 15.800 22.600 16.200 ;
        RECT 23.000 15.800 23.400 16.200 ;
        RECT 25.400 15.800 25.800 16.200 ;
        RECT 23.000 15.200 23.300 15.800 ;
        RECT 23.000 14.800 23.400 15.200 ;
        RECT 23.800 15.100 24.200 15.200 ;
        RECT 24.600 15.100 25.000 15.200 ;
        RECT 23.800 14.800 25.000 15.100 ;
        RECT 28.600 14.800 29.000 15.200 ;
        RECT 19.800 12.800 20.200 13.200 ;
        RECT 21.400 12.800 21.800 13.200 ;
        RECT 18.200 11.800 19.300 12.100 ;
        RECT 15.000 7.200 15.300 11.800 ;
        RECT 16.600 10.200 16.900 11.800 ;
        RECT 16.600 9.800 17.000 10.200 ;
        RECT 18.200 9.200 18.500 11.800 ;
        RECT 23.800 10.800 24.200 11.200 ;
        RECT 23.800 9.200 24.100 10.800 ;
        RECT 28.600 9.200 28.900 14.800 ;
        RECT 29.400 14.200 29.700 21.800 ;
        RECT 31.000 19.200 31.300 22.800 ;
        RECT 33.400 22.200 33.700 25.800 ;
        RECT 33.400 21.800 33.800 22.200 ;
        RECT 31.000 18.800 31.400 19.200 ;
        RECT 32.600 16.800 33.000 17.200 ;
        RECT 32.600 16.200 32.900 16.800 ;
        RECT 34.200 16.200 34.500 31.800 ;
        RECT 36.600 30.200 36.900 32.800 ;
        RECT 36.600 29.800 37.000 30.200 ;
        RECT 35.000 28.800 35.400 29.200 ;
        RECT 35.000 28.200 35.300 28.800 ;
        RECT 35.000 27.800 35.400 28.200 ;
        RECT 36.600 27.200 36.900 29.800 ;
        RECT 37.400 27.200 37.700 34.800 ;
        RECT 38.200 33.800 38.600 34.200 ;
        RECT 40.600 33.800 41.000 34.200 ;
        RECT 38.200 33.200 38.500 33.800 ;
        RECT 40.600 33.200 40.900 33.800 ;
        RECT 38.200 32.800 38.600 33.200 ;
        RECT 39.800 32.800 40.200 33.200 ;
        RECT 40.600 32.800 41.000 33.200 ;
        RECT 39.800 32.200 40.100 32.800 ;
        RECT 38.200 31.800 38.600 32.200 ;
        RECT 39.800 31.800 40.200 32.200 ;
        RECT 38.200 27.200 38.500 31.800 ;
        RECT 40.600 31.100 40.900 32.800 ;
        RECT 39.800 30.800 40.900 31.100 ;
        RECT 39.800 28.200 40.100 30.800 ;
        RECT 39.800 27.800 40.200 28.200 ;
        RECT 36.600 26.800 37.000 27.200 ;
        RECT 37.400 26.800 37.800 27.200 ;
        RECT 38.200 26.800 38.600 27.200 ;
        RECT 39.000 26.800 39.400 27.200 ;
        RECT 35.000 24.800 35.400 25.200 ;
        RECT 35.000 19.200 35.300 24.800 ;
        RECT 36.600 21.800 37.000 22.200 ;
        RECT 35.000 18.800 35.400 19.200 ;
        RECT 36.600 16.200 36.900 21.800 ;
        RECT 38.200 21.100 38.500 26.800 ;
        RECT 39.000 26.200 39.300 26.800 ;
        RECT 39.800 26.200 40.100 27.800 ;
        RECT 39.000 25.800 39.400 26.200 ;
        RECT 39.800 25.800 40.200 26.200 ;
        RECT 41.400 25.800 41.800 26.200 ;
        RECT 37.400 20.800 38.500 21.100 ;
        RECT 32.600 15.800 33.000 16.200 ;
        RECT 34.200 15.800 34.600 16.200 ;
        RECT 36.600 15.800 37.000 16.200 ;
        RECT 31.800 15.100 32.200 15.200 ;
        RECT 32.600 15.100 33.000 15.200 ;
        RECT 31.800 14.800 33.000 15.100 ;
        RECT 29.400 13.800 29.800 14.200 ;
        RECT 31.000 13.800 31.400 14.200 ;
        RECT 31.800 13.800 32.200 14.200 ;
        RECT 35.800 13.800 36.200 14.200 ;
        RECT 31.000 13.200 31.300 13.800 ;
        RECT 31.000 12.800 31.400 13.200 ;
        RECT 31.800 12.200 32.100 13.800 ;
        RECT 35.800 13.200 36.100 13.800 ;
        RECT 35.800 12.800 36.200 13.200 ;
        RECT 31.800 12.100 32.200 12.200 ;
        RECT 31.000 11.800 32.200 12.100 ;
        RECT 31.000 9.200 31.300 11.800 ;
        RECT 37.400 10.200 37.700 20.800 ;
        RECT 38.200 16.100 38.600 16.200 ;
        RECT 39.000 16.100 39.400 16.200 ;
        RECT 38.200 15.800 39.400 16.100 ;
        RECT 38.200 14.800 38.600 15.200 ;
        RECT 39.000 14.800 39.400 15.200 ;
        RECT 38.200 12.200 38.500 14.800 ;
        RECT 39.000 14.200 39.300 14.800 ;
        RECT 39.000 13.800 39.400 14.200 ;
        RECT 38.200 11.800 38.600 12.200 ;
        RECT 39.800 11.200 40.100 25.800 ;
        RECT 41.400 24.200 41.700 25.800 ;
        RECT 41.400 24.100 41.800 24.200 ;
        RECT 42.200 24.100 42.500 35.800 ;
        RECT 43.000 34.200 43.300 37.800 ;
        RECT 44.600 36.100 45.000 36.200 ;
        RECT 45.400 36.100 45.800 36.200 ;
        RECT 44.600 35.800 45.800 36.100 ;
        RECT 48.600 34.800 49.000 35.200 ;
        RECT 48.600 34.200 48.900 34.800 ;
        RECT 43.000 33.800 43.400 34.200 ;
        RECT 47.000 33.800 47.400 34.200 ;
        RECT 48.600 33.800 49.000 34.200 ;
        RECT 45.400 32.800 45.800 33.200 ;
        RECT 45.400 32.200 45.700 32.800 ;
        RECT 47.000 32.200 47.300 33.800 ;
        RECT 45.400 31.800 45.800 32.200 ;
        RECT 47.000 31.800 47.400 32.200 ;
        RECT 49.400 30.200 49.700 45.800 ;
        RECT 53.400 45.200 53.700 51.800 ;
        RECT 57.400 48.200 57.700 53.800 ;
        RECT 59.800 51.200 60.100 54.800 ;
        RECT 61.400 52.200 61.700 63.800 ;
        RECT 71.000 62.800 71.400 63.200 ;
        RECT 71.000 62.200 71.300 62.800 ;
        RECT 74.200 62.200 74.500 64.800 ;
        RECT 75.800 63.200 76.100 66.800 ;
        RECT 80.600 65.800 81.000 66.200 ;
        RECT 80.600 65.200 80.900 65.800 ;
        RECT 80.600 64.800 81.000 65.200 ;
        RECT 75.800 62.800 76.200 63.200 ;
        RECT 71.000 61.800 71.400 62.200 ;
        RECT 74.200 62.100 74.600 62.200 ;
        RECT 73.400 61.800 74.600 62.100 ;
        RECT 75.800 61.800 76.200 62.200 ;
        RECT 80.600 61.800 81.000 62.200 ;
        RECT 82.200 61.800 82.600 62.200 ;
        RECT 67.000 59.800 67.400 60.200 ;
        RECT 64.600 56.800 65.000 57.200 ;
        RECT 64.600 56.200 64.900 56.800 ;
        RECT 62.200 56.100 62.600 56.200 ;
        RECT 63.000 56.100 63.400 56.200 ;
        RECT 62.200 55.800 63.400 56.100 ;
        RECT 64.600 55.800 65.000 56.200 ;
        RECT 63.800 54.800 64.200 55.200 ;
        RECT 66.200 54.800 66.600 55.200 ;
        RECT 62.200 52.800 62.600 53.200 ;
        RECT 62.200 52.200 62.500 52.800 ;
        RECT 61.400 51.800 61.800 52.200 ;
        RECT 62.200 51.800 62.600 52.200 ;
        RECT 63.000 51.800 63.400 52.200 ;
        RECT 59.800 50.800 60.200 51.200 ;
        RECT 57.400 47.800 57.800 48.200 ;
        RECT 57.400 47.200 57.700 47.800 ;
        RECT 57.400 46.800 57.800 47.200 ;
        RECT 54.200 45.800 54.600 46.200 ;
        RECT 53.400 44.800 53.800 45.200 ;
        RECT 54.200 36.200 54.500 45.800 ;
        RECT 62.200 43.800 62.600 44.200 ;
        RECT 56.600 41.800 57.000 42.200 ;
        RECT 59.800 41.800 60.200 42.200 ;
        RECT 56.600 39.200 56.900 41.800 ;
        RECT 59.800 39.200 60.100 41.800 ;
        RECT 62.200 41.200 62.500 43.800 ;
        RECT 62.200 40.800 62.600 41.200 ;
        RECT 56.600 38.800 57.000 39.200 ;
        RECT 59.800 38.800 60.200 39.200 ;
        RECT 55.800 37.800 56.200 38.200 ;
        RECT 56.600 37.800 57.000 38.200 ;
        RECT 55.800 37.200 56.100 37.800 ;
        RECT 55.800 36.800 56.200 37.200 ;
        RECT 54.200 35.800 54.600 36.200 ;
        RECT 50.200 34.800 50.600 35.200 ;
        RECT 53.400 35.100 53.800 35.200 ;
        RECT 54.200 35.100 54.600 35.200 ;
        RECT 53.400 34.800 54.600 35.100 ;
        RECT 55.000 35.100 55.400 35.200 ;
        RECT 55.800 35.100 56.200 35.200 ;
        RECT 55.000 34.800 56.200 35.100 ;
        RECT 50.200 33.200 50.500 34.800 ;
        RECT 56.600 34.200 56.900 37.800 ;
        RECT 57.400 35.800 57.800 36.200 ;
        RECT 57.400 34.200 57.700 35.800 ;
        RECT 59.000 34.800 59.400 35.200 ;
        RECT 59.800 35.100 60.200 35.200 ;
        RECT 60.600 35.100 61.000 35.200 ;
        RECT 59.800 34.800 61.000 35.100 ;
        RECT 59.000 34.200 59.300 34.800 ;
        RECT 51.000 33.800 51.400 34.200 ;
        RECT 51.800 33.800 52.200 34.200 ;
        RECT 56.600 33.800 57.000 34.200 ;
        RECT 57.400 33.800 57.800 34.200 ;
        RECT 59.000 33.800 59.400 34.200 ;
        RECT 50.200 32.800 50.600 33.200 ;
        RECT 50.200 31.200 50.500 32.800 ;
        RECT 50.200 30.800 50.600 31.200 ;
        RECT 49.400 29.800 49.800 30.200 ;
        RECT 49.400 29.200 49.700 29.800 ;
        RECT 44.600 28.800 45.000 29.200 ;
        RECT 49.400 28.800 49.800 29.200 ;
        RECT 44.600 28.200 44.900 28.800 ;
        RECT 51.000 28.200 51.300 33.800 ;
        RECT 51.800 33.200 52.100 33.800 ;
        RECT 59.800 33.200 60.100 34.800 ;
        RECT 62.200 34.200 62.500 40.800 ;
        RECT 63.000 36.200 63.300 51.800 ;
        RECT 63.800 49.200 64.100 54.800 ;
        RECT 66.200 54.200 66.500 54.800 ;
        RECT 67.000 54.200 67.300 59.800 ;
        RECT 67.800 55.800 68.200 56.200 ;
        RECT 67.800 55.200 68.100 55.800 ;
        RECT 67.800 54.800 68.200 55.200 ;
        RECT 69.400 55.100 69.800 55.200 ;
        RECT 70.200 55.100 70.600 55.200 ;
        RECT 69.400 54.800 70.600 55.100 ;
        RECT 71.000 54.200 71.300 61.800 ;
        RECT 73.400 59.200 73.700 61.800 ;
        RECT 73.400 58.800 73.800 59.200 ;
        RECT 71.800 56.800 72.200 57.200 ;
        RECT 71.800 56.200 72.100 56.800 ;
        RECT 71.800 55.800 72.200 56.200 ;
        RECT 72.600 54.800 73.000 55.200 ;
        RECT 73.400 54.800 73.800 55.200 ;
        RECT 75.000 54.800 75.400 55.200 ;
        RECT 66.200 53.800 66.600 54.200 ;
        RECT 67.000 53.800 67.400 54.200 ;
        RECT 68.600 54.100 69.000 54.200 ;
        RECT 69.400 54.100 69.800 54.200 ;
        RECT 68.600 53.800 69.800 54.100 ;
        RECT 71.000 54.100 71.400 54.200 ;
        RECT 71.800 54.100 72.200 54.200 ;
        RECT 71.000 53.800 72.200 54.100 ;
        RECT 64.600 53.100 65.000 53.200 ;
        RECT 65.400 53.100 65.800 53.200 ;
        RECT 64.600 52.800 65.800 53.100 ;
        RECT 70.200 51.800 70.600 52.200 ;
        RECT 63.800 48.800 64.200 49.200 ;
        RECT 65.400 48.800 65.800 49.200 ;
        RECT 65.400 47.200 65.700 48.800 ;
        RECT 70.200 47.200 70.500 51.800 ;
        RECT 72.600 47.200 72.900 54.800 ;
        RECT 73.400 52.200 73.700 54.800 ;
        RECT 75.000 54.200 75.300 54.800 ;
        RECT 75.800 54.200 76.100 61.800 ;
        RECT 80.600 59.200 80.900 61.800 ;
        RECT 80.600 58.800 81.000 59.200 ;
        RECT 82.200 58.200 82.500 61.800 ;
        RECT 82.200 57.800 82.600 58.200 ;
        RECT 82.200 56.800 82.600 57.200 ;
        RECT 81.400 55.800 81.800 56.200 ;
        RECT 81.400 55.200 81.700 55.800 ;
        RECT 82.200 55.200 82.500 56.800 ;
        RECT 83.000 55.800 83.400 56.200 ;
        RECT 80.600 54.800 81.000 55.200 ;
        RECT 81.400 54.800 81.800 55.200 ;
        RECT 82.200 54.800 82.600 55.200 ;
        RECT 80.600 54.200 80.900 54.800 ;
        RECT 74.200 53.800 74.600 54.200 ;
        RECT 75.000 53.800 75.400 54.200 ;
        RECT 75.800 53.800 76.200 54.200 ;
        RECT 77.400 54.100 77.800 54.200 ;
        RECT 78.200 54.100 78.600 54.200 ;
        RECT 77.400 53.800 78.600 54.100 ;
        RECT 79.000 54.100 79.400 54.200 ;
        RECT 79.800 54.100 80.200 54.200 ;
        RECT 79.000 53.800 80.200 54.100 ;
        RECT 80.600 53.800 81.000 54.200 ;
        RECT 82.200 53.800 82.600 54.200 ;
        RECT 74.200 52.200 74.500 53.800 ;
        RECT 73.400 51.800 73.800 52.200 ;
        RECT 74.200 51.800 74.600 52.200 ;
        RECT 73.400 48.800 73.800 49.200 ;
        RECT 65.400 46.800 65.800 47.200 ;
        RECT 70.200 46.800 70.600 47.200 ;
        RECT 72.600 46.800 73.000 47.200 ;
        RECT 63.800 45.800 64.200 46.200 ;
        RECT 66.200 45.800 66.600 46.200 ;
        RECT 67.000 46.100 67.400 46.200 ;
        RECT 67.800 46.100 68.200 46.200 ;
        RECT 67.000 45.800 68.200 46.100 ;
        RECT 71.800 45.800 72.200 46.200 ;
        RECT 72.600 45.800 73.000 46.200 ;
        RECT 63.800 45.200 64.100 45.800 ;
        RECT 63.800 44.800 64.200 45.200 ;
        RECT 66.200 36.200 66.500 45.800 ;
        RECT 71.000 44.800 71.400 45.200 ;
        RECT 69.400 41.800 69.800 42.200 ;
        RECT 69.400 38.200 69.700 41.800 ;
        RECT 69.400 37.800 69.800 38.200 ;
        RECT 67.000 36.800 67.400 37.200 ;
        RECT 63.000 35.800 63.400 36.200 ;
        RECT 66.200 35.800 66.600 36.200 ;
        RECT 67.000 35.200 67.300 36.800 ;
        RECT 69.400 35.200 69.700 37.800 ;
        RECT 71.000 35.200 71.300 44.800 ;
        RECT 71.800 41.200 72.100 45.800 ;
        RECT 72.600 45.200 72.900 45.800 ;
        RECT 72.600 44.800 73.000 45.200 ;
        RECT 71.800 40.800 72.200 41.200 ;
        RECT 71.800 36.200 72.100 40.800 ;
        RECT 71.800 35.800 72.200 36.200 ;
        RECT 64.600 34.800 65.000 35.200 ;
        RECT 65.400 34.800 65.800 35.200 ;
        RECT 67.000 34.800 67.400 35.200 ;
        RECT 67.800 35.100 68.200 35.200 ;
        RECT 68.600 35.100 69.000 35.200 ;
        RECT 67.800 34.800 69.000 35.100 ;
        RECT 69.400 34.800 69.800 35.200 ;
        RECT 71.000 34.800 71.400 35.200 ;
        RECT 62.200 33.800 62.600 34.200 ;
        RECT 51.800 32.800 52.200 33.200 ;
        RECT 53.400 33.100 53.800 33.200 ;
        RECT 54.200 33.100 54.600 33.200 ;
        RECT 53.400 32.800 54.600 33.100 ;
        RECT 59.800 32.800 60.200 33.200 ;
        RECT 64.600 32.200 64.900 34.800 ;
        RECT 58.200 32.100 58.600 32.200 ;
        RECT 59.000 32.100 59.400 32.200 ;
        RECT 58.200 31.800 59.400 32.100 ;
        RECT 64.600 31.800 65.000 32.200 ;
        RECT 51.800 28.800 52.200 29.200 ;
        RECT 51.800 28.200 52.100 28.800 ;
        RECT 43.000 27.800 43.400 28.200 ;
        RECT 44.600 27.800 45.000 28.200 ;
        RECT 50.200 28.100 50.600 28.200 ;
        RECT 51.000 28.100 51.400 28.200 ;
        RECT 50.200 27.800 51.400 28.100 ;
        RECT 51.800 27.800 52.200 28.200 ;
        RECT 43.000 27.200 43.300 27.800 ;
        RECT 43.000 26.800 43.400 27.200 ;
        RECT 45.400 26.800 45.800 27.200 ;
        RECT 49.400 26.800 49.800 27.200 ;
        RECT 55.800 27.100 56.200 27.200 ;
        RECT 56.600 27.100 57.000 27.200 ;
        RECT 55.800 26.800 57.000 27.100 ;
        RECT 57.400 27.100 57.800 27.200 ;
        RECT 58.200 27.100 58.600 27.200 ;
        RECT 57.400 26.800 58.600 27.100 ;
        RECT 45.400 25.200 45.700 26.800 ;
        RECT 46.200 26.100 46.600 26.200 ;
        RECT 47.800 26.100 48.200 26.200 ;
        RECT 48.600 26.100 49.000 26.200 ;
        RECT 46.200 25.800 49.000 26.100 ;
        RECT 49.400 25.200 49.700 26.800 ;
        RECT 54.200 26.100 54.600 26.200 ;
        RECT 55.000 26.100 55.400 26.200 ;
        RECT 54.200 25.800 55.400 26.100 ;
        RECT 56.600 25.800 57.000 26.200 ;
        RECT 59.000 26.100 59.300 31.800 ;
        RECT 59.800 30.800 60.200 31.200 ;
        RECT 59.800 28.200 60.100 30.800 ;
        RECT 59.800 27.800 60.200 28.200 ;
        RECT 63.000 28.100 63.400 28.200 ;
        RECT 63.800 28.100 64.200 28.200 ;
        RECT 63.000 27.800 64.200 28.100 ;
        RECT 63.800 27.200 64.100 27.800 ;
        RECT 65.400 27.200 65.700 34.800 ;
        RECT 69.400 34.200 69.700 34.800 ;
        RECT 67.000 33.800 67.400 34.200 ;
        RECT 67.800 34.100 68.200 34.200 ;
        RECT 68.600 34.100 69.000 34.200 ;
        RECT 67.800 33.800 69.000 34.100 ;
        RECT 69.400 33.800 69.800 34.200 ;
        RECT 71.800 34.100 72.200 34.200 ;
        RECT 72.600 34.100 73.000 34.200 ;
        RECT 71.800 33.800 73.000 34.100 ;
        RECT 67.000 33.200 67.300 33.800 ;
        RECT 67.000 32.800 67.400 33.200 ;
        RECT 67.800 33.100 68.200 33.200 ;
        RECT 68.600 33.100 69.000 33.200 ;
        RECT 67.800 32.800 69.000 33.100 ;
        RECT 72.600 29.100 73.000 29.200 ;
        RECT 73.400 29.100 73.700 48.800 ;
        RECT 75.000 47.100 75.300 53.800 ;
        RECT 82.200 53.200 82.500 53.800 ;
        RECT 77.400 52.800 77.800 53.200 ;
        RECT 78.200 52.800 78.600 53.200 ;
        RECT 81.400 52.800 81.800 53.200 ;
        RECT 82.200 52.800 82.600 53.200 ;
        RECT 77.400 49.200 77.700 52.800 ;
        RECT 78.200 52.200 78.500 52.800 ;
        RECT 78.200 51.800 78.600 52.200 ;
        RECT 79.000 51.800 79.400 52.200 ;
        RECT 77.400 48.800 77.800 49.200 ;
        RECT 77.400 48.100 77.800 48.200 ;
        RECT 78.200 48.100 78.600 48.200 ;
        RECT 77.400 47.800 78.600 48.100 ;
        RECT 75.000 46.800 76.100 47.100 ;
        RECT 74.200 46.100 74.600 46.200 ;
        RECT 75.000 46.100 75.400 46.200 ;
        RECT 74.200 45.800 75.400 46.100 ;
        RECT 75.800 45.200 76.100 46.800 ;
        RECT 79.000 46.200 79.300 51.800 ;
        RECT 81.400 49.200 81.700 52.800 ;
        RECT 83.000 49.200 83.300 55.800 ;
        RECT 84.600 54.800 85.000 55.200 ;
        RECT 84.600 53.200 84.900 54.800 ;
        RECT 84.600 52.800 85.000 53.200 ;
        RECT 81.400 48.800 81.800 49.200 ;
        RECT 82.200 48.800 82.600 49.200 ;
        RECT 83.000 48.800 83.400 49.200 ;
        RECT 84.600 49.100 85.000 49.200 ;
        RECT 85.400 49.100 85.800 49.200 ;
        RECT 84.600 48.800 85.800 49.100 ;
        RECT 82.200 48.200 82.500 48.800 ;
        RECT 79.800 47.800 80.200 48.200 ;
        RECT 82.200 47.800 82.600 48.200 ;
        RECT 79.800 47.200 80.100 47.800 ;
        RECT 79.800 46.800 80.200 47.200 ;
        RECT 84.600 46.800 85.000 47.200 ;
        RECT 85.400 46.800 85.800 47.200 ;
        RECT 86.200 47.100 86.600 47.200 ;
        RECT 87.000 47.100 87.400 47.200 ;
        RECT 86.200 46.800 87.400 47.100 ;
        RECT 84.600 46.200 84.900 46.800 ;
        RECT 78.200 45.800 78.600 46.200 ;
        RECT 79.000 45.800 79.400 46.200 ;
        RECT 81.400 45.800 81.800 46.200 ;
        RECT 84.600 45.800 85.000 46.200 ;
        RECT 75.800 44.800 76.200 45.200 ;
        RECT 77.400 44.800 77.800 45.200 ;
        RECT 77.400 44.200 77.700 44.800 ;
        RECT 78.200 44.200 78.500 45.800 ;
        RECT 81.400 45.200 81.700 45.800 ;
        RECT 79.000 44.800 79.400 45.200 ;
        RECT 81.400 44.800 81.800 45.200 ;
        RECT 74.200 43.800 74.600 44.200 ;
        RECT 75.000 43.800 75.400 44.200 ;
        RECT 77.400 43.800 77.800 44.200 ;
        RECT 78.200 43.800 78.600 44.200 ;
        RECT 74.200 42.200 74.500 43.800 ;
        RECT 75.000 43.200 75.300 43.800 ;
        RECT 79.000 43.200 79.300 44.800 ;
        RECT 75.000 42.800 75.400 43.200 ;
        RECT 77.400 42.800 77.800 43.200 ;
        RECT 79.000 42.800 79.400 43.200 ;
        RECT 74.200 41.800 74.600 42.200 ;
        RECT 75.800 41.800 76.200 42.200 ;
        RECT 75.800 37.200 76.100 41.800 ;
        RECT 74.200 36.800 74.600 37.200 ;
        RECT 75.800 36.800 76.200 37.200 ;
        RECT 74.200 36.200 74.500 36.800 ;
        RECT 77.400 36.200 77.700 42.800 ;
        RECT 82.200 41.800 82.600 42.200 ;
        RECT 82.200 40.200 82.500 41.800 ;
        RECT 82.200 39.800 82.600 40.200 ;
        RECT 83.800 39.800 84.200 40.200 ;
        RECT 81.400 37.800 81.800 38.200 ;
        RECT 79.800 37.100 80.200 37.200 ;
        RECT 80.600 37.100 81.000 37.200 ;
        RECT 79.800 36.800 81.000 37.100 ;
        RECT 74.200 35.800 74.600 36.200 ;
        RECT 77.400 35.800 77.800 36.200 ;
        RECT 74.200 34.800 74.600 35.200 ;
        RECT 75.800 35.100 76.200 35.200 ;
        RECT 76.600 35.100 77.000 35.200 ;
        RECT 75.800 34.800 77.000 35.100 ;
        RECT 74.200 34.200 74.500 34.800 ;
        RECT 74.200 33.800 74.600 34.200 ;
        RECT 77.400 32.200 77.700 35.800 ;
        RECT 79.000 34.800 79.400 35.200 ;
        RECT 79.000 34.200 79.300 34.800 ;
        RECT 81.400 34.200 81.700 37.800 ;
        RECT 82.200 36.800 82.600 37.200 ;
        RECT 82.200 36.200 82.500 36.800 ;
        RECT 83.800 36.200 84.100 39.800 ;
        RECT 84.600 38.200 84.900 45.800 ;
        RECT 85.400 45.200 85.700 46.800 ;
        RECT 85.400 44.800 85.800 45.200 ;
        RECT 84.600 37.800 85.000 38.200 ;
        RECT 82.200 35.800 82.600 36.200 ;
        RECT 83.800 35.800 84.200 36.200 ;
        RECT 85.400 35.200 85.700 44.800 ;
        RECT 82.200 34.800 82.600 35.200 ;
        RECT 84.600 34.800 85.000 35.200 ;
        RECT 85.400 34.800 85.800 35.200 ;
        RECT 79.000 33.800 79.400 34.200 ;
        RECT 79.800 34.100 80.200 34.200 ;
        RECT 80.600 34.100 81.000 34.200 ;
        RECT 79.800 33.800 81.000 34.100 ;
        RECT 81.400 33.800 81.800 34.200 ;
        RECT 77.400 31.800 77.800 32.200 ;
        RECT 72.600 28.800 73.700 29.100 ;
        RECT 77.400 29.800 77.800 30.200 ;
        RECT 77.400 29.200 77.700 29.800 ;
        RECT 77.400 28.800 77.800 29.200 ;
        RECT 68.600 27.800 69.000 28.200 ;
        RECT 69.400 27.800 69.800 28.200 ;
        RECT 73.400 28.100 73.800 28.200 ;
        RECT 74.200 28.100 74.600 28.200 ;
        RECT 73.400 27.800 74.600 28.100 ;
        RECT 79.000 27.800 79.400 28.200 ;
        RECT 81.400 27.800 81.800 28.200 ;
        RECT 68.600 27.200 68.900 27.800 ;
        RECT 63.800 26.800 64.200 27.200 ;
        RECT 64.600 26.800 65.000 27.200 ;
        RECT 65.400 26.800 65.800 27.200 ;
        RECT 68.600 26.800 69.000 27.200 ;
        RECT 64.600 26.200 64.900 26.800 ;
        RECT 69.400 26.200 69.700 27.800 ;
        RECT 71.000 26.800 71.400 27.200 ;
        RECT 72.600 27.100 73.000 27.200 ;
        RECT 73.400 27.100 73.800 27.200 ;
        RECT 75.800 27.100 76.200 27.200 ;
        RECT 76.600 27.100 77.000 27.200 ;
        RECT 72.600 26.800 74.500 27.100 ;
        RECT 75.800 26.800 77.000 27.100 ;
        RECT 71.000 26.200 71.300 26.800 ;
        RECT 58.200 25.800 59.300 26.100 ;
        RECT 61.400 25.800 61.800 26.200 ;
        RECT 63.800 25.800 64.200 26.200 ;
        RECT 64.600 25.800 65.000 26.200 ;
        RECT 66.200 25.800 66.600 26.200 ;
        RECT 69.400 25.800 69.800 26.200 ;
        RECT 71.000 25.800 71.400 26.200 ;
        RECT 45.400 24.800 45.800 25.200 ;
        RECT 47.800 24.800 48.200 25.200 ;
        RECT 49.400 24.800 49.800 25.200 ;
        RECT 41.400 23.800 42.500 24.100 ;
        RECT 47.800 24.200 48.100 24.800 ;
        RECT 47.800 23.800 48.200 24.200 ;
        RECT 51.000 24.100 51.400 24.200 ;
        RECT 51.800 24.100 52.200 24.200 ;
        RECT 51.000 23.800 52.200 24.100 ;
        RECT 44.600 21.800 45.000 22.200 ;
        RECT 46.200 21.800 46.600 22.200 ;
        RECT 51.000 21.800 51.400 22.200 ;
        RECT 52.600 21.800 53.000 22.200 ;
        RECT 55.800 21.800 56.200 22.200 ;
        RECT 44.600 20.200 44.900 21.800 ;
        RECT 44.600 19.800 45.000 20.200 ;
        RECT 45.400 16.800 45.800 17.200 ;
        RECT 44.600 15.800 45.000 16.200 ;
        RECT 40.600 15.100 41.000 15.200 ;
        RECT 41.400 15.100 41.800 15.200 ;
        RECT 40.600 14.800 41.800 15.100 ;
        RECT 41.400 13.800 41.800 14.200 ;
        RECT 43.800 14.000 44.200 14.400 ;
        RECT 44.600 14.200 44.900 15.800 ;
        RECT 45.400 15.200 45.700 16.800 ;
        RECT 46.200 16.200 46.500 21.800 ;
        RECT 46.200 15.800 46.600 16.200 ;
        RECT 47.800 15.800 48.200 16.200 ;
        RECT 45.400 14.800 45.800 15.200 ;
        RECT 47.800 14.200 48.100 15.800 ;
        RECT 48.600 14.800 49.000 15.200 ;
        RECT 49.400 15.100 49.800 15.200 ;
        RECT 50.200 15.100 50.600 15.200 ;
        RECT 49.400 14.800 50.600 15.100 ;
        RECT 41.400 11.200 41.700 13.800 ;
        RECT 43.800 13.200 44.100 14.000 ;
        RECT 44.600 13.800 45.000 14.200 ;
        RECT 45.400 13.800 45.800 14.200 ;
        RECT 47.800 13.800 48.200 14.200 ;
        RECT 45.400 13.200 45.700 13.800 ;
        RECT 43.800 12.800 44.200 13.200 ;
        RECT 45.400 12.800 45.800 13.200 ;
        RECT 47.000 13.100 47.400 13.200 ;
        RECT 47.800 13.100 48.200 13.200 ;
        RECT 47.000 12.800 48.200 13.100 ;
        RECT 48.600 12.200 48.900 14.800 ;
        RECT 51.000 14.200 51.300 21.800 ;
        RECT 52.600 16.200 52.900 21.800 ;
        RECT 55.800 19.200 56.100 21.800 ;
        RECT 55.800 18.800 56.200 19.200 ;
        RECT 54.200 17.800 54.600 18.200 ;
        RECT 52.600 15.800 53.000 16.200 ;
        RECT 53.400 15.800 53.800 16.200 ;
        RECT 53.400 15.200 53.700 15.800 ;
        RECT 51.800 14.800 52.200 15.200 ;
        RECT 53.400 14.800 53.800 15.200 ;
        RECT 49.400 13.800 49.800 14.200 ;
        RECT 51.000 13.800 51.400 14.200 ;
        RECT 49.400 13.200 49.700 13.800 ;
        RECT 49.400 12.800 49.800 13.200 ;
        RECT 42.200 11.800 42.600 12.200 ;
        RECT 48.600 11.800 49.000 12.200 ;
        RECT 39.800 10.800 40.200 11.200 ;
        RECT 41.400 10.800 41.800 11.200 ;
        RECT 34.200 9.800 34.600 10.200 ;
        RECT 37.400 9.800 37.800 10.200 ;
        RECT 34.200 9.200 34.500 9.800 ;
        RECT 18.200 8.800 18.600 9.200 ;
        RECT 23.800 8.800 24.200 9.200 ;
        RECT 28.600 8.800 29.000 9.200 ;
        RECT 31.000 8.800 31.400 9.200 ;
        RECT 34.200 8.800 34.600 9.200 ;
        RECT 41.400 8.800 41.800 9.200 ;
        RECT 41.400 8.200 41.700 8.800 ;
        RECT 15.700 7.500 16.100 7.900 ;
        RECT 19.000 7.500 19.400 7.900 ;
        RECT 5.000 6.700 5.400 6.800 ;
        RECT 7.100 5.100 7.400 6.800 ;
        RECT 13.400 6.600 13.800 7.000 ;
        RECT 14.200 6.800 14.600 7.200 ;
        RECT 15.000 6.800 15.400 7.200 ;
        RECT 10.200 6.100 10.600 6.200 ;
        RECT 11.000 6.100 11.400 6.200 ;
        RECT 10.200 5.800 11.400 6.100 ;
        RECT 3.700 4.700 4.100 5.100 ;
        RECT 7.000 4.700 7.400 5.100 ;
        RECT 15.700 5.100 16.000 7.500 ;
        RECT 19.100 7.100 19.400 7.500 ;
        RECT 17.000 6.800 19.400 7.100 ;
        RECT 17.000 6.700 17.400 6.800 ;
        RECT 19.100 5.100 19.400 6.800 ;
        RECT 15.700 4.700 16.100 5.100 ;
        RECT 19.000 4.700 19.400 5.100 ;
        RECT 21.400 7.500 21.800 7.900 ;
        RECT 24.500 7.800 24.900 7.900 ;
        RECT 41.400 7.800 41.800 8.200 ;
        RECT 22.100 7.500 24.900 7.800 ;
        RECT 21.400 7.100 21.700 7.500 ;
        RECT 22.100 7.400 22.500 7.500 ;
        RECT 23.800 7.400 24.200 7.500 ;
        RECT 21.400 6.800 24.200 7.100 ;
        RECT 21.400 5.100 21.700 6.800 ;
        RECT 23.900 6.100 24.200 6.800 ;
        RECT 23.900 5.700 24.300 6.100 ;
        RECT 24.600 5.100 24.900 7.500 ;
        RECT 42.200 7.200 42.500 11.800 ;
        RECT 51.000 10.800 51.400 11.200 ;
        RECT 44.600 9.800 45.000 10.200 ;
        RECT 43.800 8.800 44.200 9.200 ;
        RECT 21.400 4.700 21.800 5.100 ;
        RECT 24.500 4.700 24.900 5.100 ;
        RECT 37.400 6.800 37.800 7.200 ;
        RECT 41.400 6.800 41.800 7.200 ;
        RECT 42.200 6.800 42.600 7.200 ;
        RECT 37.400 5.200 37.700 6.800 ;
        RECT 41.400 6.200 41.700 6.800 ;
        RECT 43.800 6.200 44.100 8.800 ;
        RECT 44.600 7.200 44.900 9.800 ;
        RECT 47.000 8.800 47.400 9.200 ;
        RECT 45.400 8.100 45.800 8.200 ;
        RECT 46.200 8.100 46.600 8.200 ;
        RECT 45.400 7.800 46.600 8.100 ;
        RECT 47.000 7.200 47.300 8.800 ;
        RECT 51.000 8.200 51.300 10.800 ;
        RECT 51.800 9.200 52.100 14.800 ;
        RECT 54.200 14.200 54.500 17.800 ;
        RECT 55.000 16.100 55.400 16.200 ;
        RECT 55.800 16.100 56.200 16.200 ;
        RECT 55.000 15.800 56.200 16.100 ;
        RECT 56.600 15.200 56.900 25.800 ;
        RECT 57.400 17.800 57.800 18.200 ;
        RECT 57.400 17.200 57.700 17.800 ;
        RECT 57.400 16.800 57.800 17.200 ;
        RECT 58.200 15.200 58.500 25.800 ;
        RECT 61.400 25.200 61.700 25.800 ;
        RECT 59.000 24.800 59.400 25.200 ;
        RECT 61.400 24.800 61.800 25.200 ;
        RECT 55.000 14.800 55.400 15.200 ;
        RECT 56.600 14.800 57.000 15.200 ;
        RECT 58.200 14.800 58.600 15.200 ;
        RECT 52.600 14.100 53.000 14.200 ;
        RECT 53.400 14.100 53.800 14.200 ;
        RECT 52.600 13.800 53.800 14.100 ;
        RECT 54.200 13.800 54.600 14.200 ;
        RECT 55.000 11.200 55.300 14.800 ;
        RECT 59.000 14.200 59.300 24.800 ;
        RECT 62.200 15.100 62.600 15.200 ;
        RECT 63.000 15.100 63.400 15.200 ;
        RECT 62.200 14.800 63.400 15.100 ;
        RECT 58.200 13.800 58.600 14.200 ;
        RECT 59.000 13.800 59.400 14.200 ;
        RECT 59.800 14.000 60.200 14.400 ;
        RECT 63.800 14.200 64.100 25.800 ;
        RECT 58.200 12.200 58.500 13.800 ;
        RECT 55.800 11.800 56.200 12.200 ;
        RECT 58.200 11.800 58.600 12.200 ;
        RECT 52.600 10.800 53.000 11.200 ;
        RECT 55.000 10.800 55.400 11.200 ;
        RECT 52.600 9.200 52.900 10.800 ;
        RECT 55.800 9.200 56.100 11.800 ;
        RECT 59.000 11.200 59.300 13.800 ;
        RECT 59.800 12.200 60.100 14.000 ;
        RECT 63.800 13.800 64.200 14.200 ;
        RECT 64.600 12.200 64.900 25.800 ;
        RECT 66.200 25.200 66.500 25.800 ;
        RECT 66.200 24.800 66.600 25.200 ;
        RECT 67.000 24.800 67.400 25.200 ;
        RECT 69.400 24.800 69.800 25.200 ;
        RECT 67.000 24.200 67.300 24.800 ;
        RECT 67.000 23.800 67.400 24.200 ;
        RECT 69.400 21.200 69.700 24.800 ;
        RECT 67.000 20.800 67.400 21.200 ;
        RECT 69.400 20.800 69.800 21.200 ;
        RECT 65.400 19.800 65.800 20.200 ;
        RECT 59.800 11.800 60.200 12.200 ;
        RECT 63.000 11.800 63.400 12.200 ;
        RECT 64.600 11.800 65.000 12.200 ;
        RECT 59.000 10.800 59.400 11.200 ;
        RECT 63.000 9.200 63.300 11.800 ;
        RECT 51.800 8.800 52.200 9.200 ;
        RECT 52.600 8.800 53.000 9.200 ;
        RECT 55.800 8.800 56.200 9.200 ;
        RECT 63.000 8.800 63.400 9.200 ;
        RECT 63.000 8.200 63.300 8.800 ;
        RECT 51.000 7.800 51.400 8.200 ;
        RECT 60.600 7.800 61.000 8.200 ;
        RECT 63.000 7.800 63.400 8.200 ;
        RECT 51.000 7.200 51.300 7.800 ;
        RECT 60.600 7.200 60.900 7.800 ;
        RECT 65.400 7.200 65.700 19.800 ;
        RECT 66.200 15.800 66.600 16.200 ;
        RECT 66.200 15.200 66.500 15.800 ;
        RECT 67.000 15.200 67.300 20.800 ;
        RECT 71.800 18.800 72.200 19.200 ;
        RECT 68.600 15.800 69.000 16.200 ;
        RECT 68.600 15.200 68.900 15.800 ;
        RECT 66.200 14.800 66.600 15.200 ;
        RECT 67.000 14.800 67.400 15.200 ;
        RECT 68.600 14.800 69.000 15.200 ;
        RECT 70.200 15.100 70.600 15.200 ;
        RECT 71.000 15.100 71.400 15.200 ;
        RECT 70.200 14.800 71.400 15.100 ;
        RECT 71.800 14.200 72.100 18.800 ;
        RECT 74.200 15.200 74.500 26.800 ;
        RECT 79.000 15.200 79.300 27.800 ;
        RECT 80.600 26.800 81.000 27.200 ;
        RECT 79.800 24.800 80.200 25.200 ;
        RECT 79.800 24.200 80.100 24.800 ;
        RECT 79.800 23.800 80.200 24.200 ;
        RECT 80.600 20.200 80.900 26.800 ;
        RECT 81.400 26.200 81.700 27.800 ;
        RECT 82.200 27.200 82.500 34.800 ;
        RECT 84.600 34.200 84.900 34.800 ;
        RECT 84.600 33.800 85.000 34.200 ;
        RECT 82.200 26.800 82.600 27.200 ;
        RECT 81.400 25.800 81.800 26.200 ;
        RECT 84.600 25.800 85.000 26.200 ;
        RECT 82.200 25.100 82.600 25.200 ;
        RECT 83.000 25.100 83.400 25.200 ;
        RECT 82.200 24.800 83.400 25.100 ;
        RECT 84.600 22.200 84.900 25.800 ;
        RECT 84.600 21.800 85.000 22.200 ;
        RECT 85.400 21.800 85.800 22.200 ;
        RECT 80.600 19.800 81.000 20.200 ;
        RECT 83.000 16.800 83.400 17.200 ;
        RECT 83.000 16.200 83.300 16.800 ;
        RECT 79.800 16.100 80.200 16.200 ;
        RECT 80.600 16.100 81.000 16.200 ;
        RECT 79.800 15.800 81.000 16.100 ;
        RECT 83.000 15.800 83.400 16.200 ;
        RECT 84.600 15.200 84.900 21.800 ;
        RECT 85.400 19.200 85.700 21.800 ;
        RECT 85.400 18.800 85.800 19.200 ;
        RECT 74.200 14.800 74.600 15.200 ;
        RECT 77.400 14.800 77.800 15.200 ;
        RECT 78.200 14.800 78.600 15.200 ;
        RECT 79.000 14.800 79.400 15.200 ;
        RECT 79.800 15.100 80.200 15.200 ;
        RECT 80.600 15.100 81.000 15.200 ;
        RECT 79.800 14.800 81.000 15.100 ;
        RECT 82.200 15.100 82.600 15.200 ;
        RECT 83.000 15.100 83.400 15.200 ;
        RECT 82.200 14.800 83.400 15.100 ;
        RECT 84.600 14.800 85.000 15.200 ;
        RECT 77.400 14.200 77.700 14.800 ;
        RECT 67.000 14.100 67.400 14.200 ;
        RECT 67.800 14.100 68.200 14.200 ;
        RECT 67.000 13.800 68.200 14.100 ;
        RECT 69.400 13.800 69.800 14.200 ;
        RECT 71.800 13.800 72.200 14.200 ;
        RECT 75.000 13.800 75.400 14.200 ;
        RECT 77.400 13.800 77.800 14.200 ;
        RECT 69.400 13.200 69.700 13.800 ;
        RECT 75.000 13.200 75.300 13.800 ;
        RECT 69.400 12.800 69.800 13.200 ;
        RECT 71.000 12.800 71.400 13.200 ;
        RECT 71.800 12.800 72.200 13.200 ;
        RECT 75.000 12.800 75.400 13.200 ;
        RECT 76.600 12.800 77.000 13.200 ;
        RECT 71.000 12.200 71.300 12.800 ;
        RECT 66.200 12.100 66.600 12.200 ;
        RECT 67.000 12.100 67.400 12.200 ;
        RECT 66.200 11.800 67.400 12.100 ;
        RECT 71.000 11.800 71.400 12.200 ;
        RECT 71.800 9.200 72.100 12.800 ;
        RECT 76.600 12.200 76.900 12.800 ;
        RECT 73.400 12.100 73.800 12.200 ;
        RECT 74.200 12.100 74.600 12.200 ;
        RECT 73.400 11.800 74.600 12.100 ;
        RECT 75.800 11.800 76.200 12.200 ;
        RECT 76.600 11.800 77.000 12.200 ;
        RECT 75.800 11.200 76.100 11.800 ;
        RECT 75.800 10.800 76.200 11.200 ;
        RECT 77.400 10.200 77.700 13.800 ;
        RECT 73.400 9.800 73.800 10.200 ;
        RECT 77.400 9.800 77.800 10.200 ;
        RECT 67.800 8.800 68.200 9.200 ;
        RECT 71.800 8.800 72.200 9.200 ;
        RECT 66.200 7.800 66.600 8.200 ;
        RECT 44.600 7.100 45.000 7.200 ;
        RECT 44.600 6.800 45.700 7.100 ;
        RECT 47.000 6.800 47.400 7.200 ;
        RECT 47.800 7.100 48.200 7.200 ;
        RECT 48.600 7.100 49.000 7.200 ;
        RECT 47.800 6.800 49.000 7.100 ;
        RECT 51.000 6.800 51.400 7.200 ;
        RECT 52.600 6.800 53.000 7.200 ;
        RECT 60.600 7.100 61.000 7.200 ;
        RECT 61.400 7.100 61.800 7.200 ;
        RECT 60.600 6.800 61.800 7.100 ;
        RECT 63.000 6.800 63.400 7.200 ;
        RECT 65.400 6.800 65.800 7.200 ;
        RECT 39.000 6.100 39.400 6.200 ;
        RECT 39.800 6.100 40.200 6.200 ;
        RECT 39.000 5.800 40.200 6.100 ;
        RECT 41.400 5.800 41.800 6.200 ;
        RECT 42.200 5.800 42.600 6.200 ;
        RECT 43.800 5.800 44.200 6.200 ;
        RECT 42.200 5.200 42.500 5.800 ;
        RECT 45.400 5.200 45.700 6.800 ;
        RECT 52.600 6.200 52.900 6.800 ;
        RECT 63.000 6.200 63.300 6.800 ;
        RECT 66.200 6.200 66.500 7.800 ;
        RECT 49.400 6.100 49.800 6.200 ;
        RECT 50.200 6.100 50.600 6.200 ;
        RECT 49.400 5.800 50.600 6.100 ;
        RECT 52.600 5.800 53.000 6.200 ;
        RECT 63.000 5.800 63.400 6.200 ;
        RECT 66.200 5.800 66.600 6.200 ;
        RECT 67.800 5.200 68.100 8.800 ;
        RECT 69.300 7.500 69.700 7.900 ;
        RECT 70.200 7.500 72.300 7.800 ;
        RECT 72.600 7.500 73.000 7.900 ;
        RECT 37.400 4.800 37.800 5.200 ;
        RECT 42.200 4.800 42.600 5.200 ;
        RECT 45.400 4.800 45.800 5.200 ;
        RECT 63.800 5.100 64.200 5.200 ;
        RECT 64.600 5.100 65.000 5.200 ;
        RECT 63.800 4.800 65.000 5.100 ;
        RECT 67.000 5.100 67.400 5.200 ;
        RECT 67.800 5.100 68.200 5.200 ;
        RECT 67.000 4.800 68.200 5.100 ;
        RECT 69.300 5.100 69.600 7.500 ;
        RECT 70.200 7.400 70.600 7.500 ;
        RECT 71.900 7.400 72.300 7.500 ;
        RECT 72.700 7.100 73.000 7.500 ;
        RECT 70.600 6.800 73.000 7.100 ;
        RECT 73.400 7.200 73.700 9.800 ;
        RECT 78.200 9.200 78.500 14.800 ;
        RECT 79.800 13.800 80.200 14.200 ;
        RECT 82.200 14.100 82.600 14.200 ;
        RECT 83.000 14.100 83.400 14.200 ;
        RECT 82.200 13.800 83.400 14.100 ;
        RECT 79.000 9.800 79.400 10.200 ;
        RECT 78.200 8.800 78.600 9.200 ;
        RECT 74.900 7.500 75.300 7.900 ;
        RECT 75.800 7.500 77.900 7.800 ;
        RECT 78.200 7.500 78.600 7.900 ;
        RECT 73.400 6.800 73.800 7.200 ;
        RECT 74.200 6.800 74.600 7.200 ;
        RECT 70.600 6.700 71.000 6.800 ;
        RECT 72.700 5.100 73.000 6.800 ;
        RECT 74.200 6.200 74.500 6.800 ;
        RECT 74.200 5.800 74.600 6.200 ;
        RECT 69.300 4.700 69.700 5.100 ;
        RECT 72.600 4.700 73.000 5.100 ;
        RECT 74.900 5.100 75.200 7.500 ;
        RECT 75.800 7.400 76.200 7.500 ;
        RECT 77.500 7.400 77.900 7.500 ;
        RECT 78.300 7.100 78.600 7.500 ;
        RECT 76.200 6.800 78.600 7.100 ;
        RECT 79.000 7.200 79.300 9.800 ;
        RECT 79.800 8.200 80.100 13.800 ;
        RECT 83.800 13.100 84.200 13.200 ;
        RECT 84.600 13.100 85.000 13.200 ;
        RECT 83.800 12.800 85.000 13.100 ;
        RECT 83.800 10.800 84.200 11.200 ;
        RECT 79.800 7.800 80.200 8.200 ;
        RECT 79.000 6.800 79.400 7.200 ;
        RECT 81.400 6.800 81.800 7.200 ;
        RECT 76.200 6.700 76.600 6.800 ;
        RECT 78.300 5.100 78.600 6.800 ;
        RECT 81.400 6.200 81.700 6.800 ;
        RECT 79.000 6.100 79.400 6.200 ;
        RECT 79.800 6.100 80.200 6.200 ;
        RECT 79.000 5.800 80.200 6.100 ;
        RECT 81.400 5.800 81.800 6.200 ;
        RECT 74.900 4.700 75.300 5.100 ;
        RECT 78.200 4.700 78.600 5.100 ;
        RECT 83.800 5.200 84.100 10.800 ;
        RECT 83.800 4.800 84.200 5.200 ;
      LAYER via2 ;
        RECT 3.000 66.800 3.400 67.200 ;
        RECT 39.000 66.800 39.400 67.200 ;
        RECT 43.800 66.800 44.200 67.200 ;
        RECT 44.600 65.800 45.000 66.200 ;
        RECT 19.800 53.800 20.200 54.200 ;
        RECT 3.000 45.800 3.400 46.200 ;
        RECT 7.000 45.800 7.400 46.200 ;
        RECT 7.000 44.800 7.400 45.200 ;
        RECT 7.000 35.800 7.400 36.200 ;
        RECT 7.000 24.800 7.400 25.200 ;
        RECT 5.400 14.800 5.800 15.200 ;
        RECT 7.000 13.800 7.400 14.200 ;
        RECT 22.200 46.800 22.600 47.200 ;
        RECT 35.800 46.800 36.200 47.200 ;
        RECT 68.600 64.800 69.000 65.200 ;
        RECT 59.000 56.800 59.400 57.200 ;
        RECT 53.400 54.800 53.800 55.200 ;
        RECT 52.600 47.800 53.000 48.200 ;
        RECT 50.200 45.800 50.600 46.200 ;
        RECT 20.600 35.800 21.000 36.200 ;
        RECT 3.000 5.800 3.400 6.200 ;
        RECT 16.600 14.800 17.000 15.200 ;
        RECT 42.200 42.800 42.600 43.200 ;
        RECT 18.200 12.800 18.600 13.200 ;
        RECT 31.800 11.800 32.200 12.200 ;
        RECT 74.200 61.800 74.600 62.200 ;
        RECT 60.600 34.800 61.000 35.200 ;
        RECT 71.800 53.800 72.200 54.200 ;
        RECT 78.200 53.800 78.600 54.200 ;
        RECT 54.200 32.800 54.600 33.200 ;
        RECT 59.000 31.800 59.400 32.200 ;
        RECT 58.200 26.800 58.600 27.200 ;
        RECT 47.800 25.800 48.200 26.200 ;
        RECT 55.000 25.800 55.400 26.200 ;
        RECT 63.800 27.800 64.200 28.200 ;
        RECT 78.200 47.800 78.600 48.200 ;
        RECT 80.600 36.800 81.000 37.200 ;
        RECT 41.400 14.800 41.800 15.200 ;
        RECT 47.800 12.800 48.200 13.200 ;
        RECT 46.200 7.800 46.600 8.200 ;
        RECT 53.400 13.800 53.800 14.200 ;
        RECT 71.000 14.800 71.400 15.200 ;
        RECT 80.600 15.800 81.000 16.200 ;
        RECT 80.600 14.800 81.000 15.200 ;
        RECT 83.000 14.800 83.400 15.200 ;
        RECT 67.000 11.800 67.400 12.200 ;
        RECT 74.200 11.800 74.600 12.200 ;
        RECT 61.400 6.800 61.800 7.200 ;
        RECT 39.800 5.800 40.200 6.200 ;
        RECT 50.200 5.800 50.600 6.200 ;
        RECT 64.600 4.800 65.000 5.200 ;
        RECT 79.800 5.800 80.200 6.200 ;
      LAYER metal3 ;
        RECT 20.600 68.100 21.000 68.200 ;
        RECT 23.800 68.100 24.200 68.200 ;
        RECT 31.800 68.100 32.200 68.200 ;
        RECT 38.200 68.100 38.600 68.200 ;
        RECT 20.600 67.800 38.600 68.100 ;
        RECT 46.200 68.100 46.600 68.200 ;
        RECT 49.400 68.100 49.800 68.200 ;
        RECT 67.000 68.100 67.400 68.200 ;
        RECT 46.200 67.800 67.400 68.100 ;
        RECT 3.000 67.100 3.400 67.200 ;
        RECT 9.400 67.100 9.800 67.200 ;
        RECT 3.000 66.800 9.800 67.100 ;
        RECT 17.400 67.100 17.800 67.200 ;
        RECT 25.400 67.100 25.800 67.200 ;
        RECT 17.400 66.800 25.800 67.100 ;
        RECT 33.400 67.100 33.800 67.200 ;
        RECT 39.000 67.100 39.400 67.200 ;
        RECT 43.800 67.100 44.200 67.200 ;
        RECT 33.400 66.800 37.700 67.100 ;
        RECT 39.000 66.800 44.200 67.100 ;
        RECT 48.600 67.100 49.000 67.200 ;
        RECT 48.600 66.800 50.500 67.100 ;
        RECT 37.400 66.200 37.700 66.800 ;
        RECT 50.200 66.200 50.500 66.800 ;
        RECT 53.400 66.800 53.800 67.200 ;
        RECT 10.200 66.100 10.600 66.200 ;
        RECT 12.600 66.100 13.000 66.200 ;
        RECT 10.200 65.800 13.000 66.100 ;
        RECT 25.400 66.100 25.800 66.200 ;
        RECT 31.000 66.100 31.400 66.200 ;
        RECT 25.400 65.800 31.400 66.100 ;
        RECT 37.400 65.800 37.800 66.200 ;
        RECT 41.400 65.800 41.800 66.200 ;
        RECT 44.600 66.100 45.000 66.200 ;
        RECT 46.200 66.100 46.600 66.200 ;
        RECT 44.600 65.800 46.600 66.100 ;
        RECT 50.200 66.100 50.600 66.200 ;
        RECT 53.400 66.100 53.700 66.800 ;
        RECT 50.200 65.800 53.700 66.100 ;
        RECT 75.000 65.800 75.400 66.200 ;
        RECT 80.600 65.800 81.000 66.200 ;
        RECT 29.400 65.100 29.800 65.200 ;
        RECT 41.400 65.100 41.700 65.800 ;
        RECT 45.400 65.100 45.800 65.200 ;
        RECT 29.400 64.800 40.900 65.100 ;
        RECT 41.400 64.800 45.800 65.100 ;
        RECT 52.600 65.100 53.000 65.200 ;
        RECT 54.200 65.100 54.600 65.200 ;
        RECT 52.600 64.800 54.600 65.100 ;
        RECT 68.600 65.100 69.000 65.200 ;
        RECT 75.000 65.100 75.300 65.800 ;
        RECT 68.600 64.800 75.300 65.100 ;
        RECT 80.600 65.200 80.900 65.800 ;
        RECT 80.600 64.800 81.000 65.200 ;
        RECT 19.000 64.100 19.400 64.200 ;
        RECT 11.000 63.800 19.400 64.100 ;
        RECT 40.600 64.100 40.900 64.800 ;
        RECT 43.800 64.100 44.200 64.200 ;
        RECT 40.600 63.800 44.200 64.100 ;
        RECT 11.000 63.200 11.300 63.800 ;
        RECT 11.000 62.800 11.400 63.200 ;
        RECT 71.000 63.100 71.400 63.200 ;
        RECT 75.800 63.100 76.200 63.200 ;
        RECT 71.000 62.800 76.200 63.100 ;
        RECT 27.000 62.100 27.400 62.200 ;
        RECT 34.200 62.100 34.600 62.200 ;
        RECT 27.000 61.800 34.600 62.100 ;
        RECT 74.200 62.100 74.600 62.200 ;
        RECT 75.800 62.100 76.200 62.200 ;
        RECT 74.200 61.800 76.200 62.100 ;
        RECT 55.800 60.100 56.200 60.200 ;
        RECT 67.000 60.100 67.400 60.200 ;
        RECT 55.800 59.800 67.400 60.100 ;
        RECT 35.000 59.100 35.400 59.200 ;
        RECT 43.800 59.100 44.200 59.200 ;
        RECT 45.400 59.100 45.800 59.200 ;
        RECT 35.000 58.800 45.800 59.100 ;
        RECT 80.600 59.100 81.000 59.200 ;
        RECT 84.600 59.100 85.000 59.200 ;
        RECT 80.600 58.800 85.000 59.100 ;
        RECT 12.600 58.100 13.000 58.200 ;
        RECT 42.200 58.100 42.600 58.200 ;
        RECT 12.600 57.800 42.600 58.100 ;
        RECT 82.200 58.100 82.600 58.200 ;
        RECT 83.000 58.100 83.400 58.200 ;
        RECT 82.200 57.800 83.400 58.100 ;
        RECT 7.800 57.100 8.200 57.200 ;
        RECT 11.000 57.100 11.400 57.200 ;
        RECT 22.200 57.100 22.600 57.200 ;
        RECT 35.800 57.100 36.200 57.200 ;
        RECT 7.800 56.800 36.200 57.100 ;
        RECT 59.000 57.100 59.400 57.200 ;
        RECT 60.600 57.100 61.000 57.200 ;
        RECT 71.800 57.100 72.200 57.200 ;
        RECT 82.200 57.100 82.600 57.200 ;
        RECT 59.000 56.800 82.600 57.100 ;
        RECT 1.400 56.100 1.800 56.200 ;
        RECT 4.600 56.100 5.000 56.200 ;
        RECT 1.400 55.800 5.000 56.100 ;
        RECT 10.200 55.800 10.600 56.200 ;
        RECT 14.200 56.100 14.600 56.200 ;
        RECT 18.200 56.100 18.600 56.200 ;
        RECT 14.200 55.800 18.600 56.100 ;
        RECT 43.000 56.100 43.400 56.200 ;
        RECT 50.200 56.100 50.600 56.200 ;
        RECT 43.000 55.800 50.600 56.100 ;
        RECT 52.600 56.100 53.000 56.200 ;
        RECT 53.400 56.100 53.800 56.200 ;
        RECT 52.600 55.800 53.800 56.100 ;
        RECT 59.800 56.100 60.200 56.200 ;
        RECT 62.200 56.100 62.600 56.200 ;
        RECT 59.800 55.800 62.600 56.100 ;
        RECT 64.600 56.100 65.000 56.200 ;
        RECT 67.800 56.100 68.200 56.200 ;
        RECT 64.600 55.800 68.200 56.100 ;
        RECT 81.400 55.800 81.800 56.200 ;
        RECT 1.400 55.100 1.800 55.200 ;
        RECT 3.000 55.100 3.400 55.200 ;
        RECT 10.200 55.100 10.500 55.800 ;
        RECT 1.400 54.800 10.500 55.100 ;
        RECT 39.000 55.100 39.400 55.200 ;
        RECT 47.000 55.100 47.400 55.200 ;
        RECT 39.000 54.800 47.400 55.100 ;
        RECT 53.400 55.100 53.800 55.200 ;
        RECT 59.000 55.100 59.400 55.200 ;
        RECT 53.400 54.800 59.400 55.100 ;
        RECT 59.800 55.100 60.200 55.200 ;
        RECT 66.200 55.100 66.600 55.200 ;
        RECT 59.800 54.800 66.600 55.100 ;
        RECT 69.400 55.100 69.800 55.200 ;
        RECT 72.600 55.100 73.000 55.200 ;
        RECT 81.400 55.100 81.700 55.800 ;
        RECT 69.400 54.800 81.700 55.100 ;
        RECT 5.400 54.100 5.800 54.200 ;
        RECT 7.800 54.100 8.200 54.200 ;
        RECT 5.400 53.800 8.200 54.100 ;
        RECT 9.400 54.100 9.800 54.200 ;
        RECT 14.200 54.100 14.600 54.200 ;
        RECT 9.400 53.800 14.600 54.100 ;
        RECT 19.800 54.100 20.200 54.200 ;
        RECT 23.000 54.100 23.400 54.200 ;
        RECT 19.800 53.800 23.400 54.100 ;
        RECT 57.400 54.100 57.800 54.200 ;
        RECT 68.600 54.100 69.000 54.200 ;
        RECT 57.400 53.800 69.000 54.100 ;
        RECT 71.800 54.100 72.200 54.200 ;
        RECT 75.000 54.100 75.400 54.200 ;
        RECT 71.800 53.800 75.400 54.100 ;
        RECT 78.200 54.100 78.600 54.200 ;
        RECT 79.000 54.100 79.400 54.200 ;
        RECT 78.200 53.800 79.400 54.100 ;
        RECT 80.600 54.100 81.000 54.200 ;
        RECT 82.200 54.100 82.600 54.200 ;
        RECT 80.600 53.800 82.600 54.100 ;
        RECT 25.400 53.100 25.800 53.200 ;
        RECT 27.000 53.100 27.400 53.200 ;
        RECT 64.600 53.100 65.000 53.200 ;
        RECT 81.400 53.100 81.800 53.200 ;
        RECT 84.600 53.100 85.000 53.200 ;
        RECT 25.400 52.800 34.500 53.100 ;
        RECT 64.600 52.800 78.500 53.100 ;
        RECT 81.400 52.800 85.000 53.100 ;
        RECT 34.200 52.100 34.500 52.800 ;
        RECT 78.200 52.200 78.500 52.800 ;
        RECT 53.400 52.100 53.800 52.200 ;
        RECT 61.400 52.100 61.800 52.200 ;
        RECT 34.200 51.800 61.800 52.100 ;
        RECT 62.200 52.100 62.600 52.200 ;
        RECT 63.000 52.100 63.400 52.200 ;
        RECT 70.200 52.100 70.600 52.200 ;
        RECT 73.400 52.100 73.800 52.200 ;
        RECT 62.200 51.800 73.800 52.100 ;
        RECT 74.200 52.100 74.600 52.200 ;
        RECT 75.000 52.100 75.400 52.200 ;
        RECT 74.200 51.800 75.400 52.100 ;
        RECT 78.200 51.800 78.600 52.200 ;
        RECT 16.600 51.100 17.000 51.200 ;
        RECT 35.800 51.100 36.200 51.200 ;
        RECT 16.600 50.800 36.200 51.100 ;
        RECT 36.600 51.100 37.000 51.200 ;
        RECT 37.400 51.100 37.800 51.200 ;
        RECT 47.000 51.100 47.400 51.200 ;
        RECT 57.400 51.100 57.800 51.200 ;
        RECT 59.800 51.100 60.200 51.200 ;
        RECT 36.600 50.800 60.200 51.100 ;
        RECT 11.800 50.100 12.200 50.200 ;
        RECT 19.000 50.100 19.400 50.200 ;
        RECT 11.800 49.800 19.400 50.100 ;
        RECT 19.800 50.100 20.200 50.200 ;
        RECT 36.600 50.100 37.000 50.200 ;
        RECT 19.800 49.800 37.000 50.100 ;
        RECT 4.600 49.100 5.000 49.200 ;
        RECT 16.600 49.100 17.000 49.200 ;
        RECT 4.600 48.800 17.000 49.100 ;
        RECT 34.200 49.100 34.600 49.200 ;
        RECT 39.800 49.100 40.200 49.200 ;
        RECT 49.400 49.100 49.800 49.200 ;
        RECT 65.400 49.100 65.800 49.200 ;
        RECT 34.200 48.800 65.800 49.100 ;
        RECT 73.400 49.100 73.800 49.200 ;
        RECT 77.400 49.100 77.800 49.200 ;
        RECT 82.200 49.100 82.600 49.200 ;
        RECT 73.400 48.800 82.600 49.100 ;
        RECT 83.000 49.100 83.400 49.200 ;
        RECT 84.600 49.100 85.000 49.200 ;
        RECT 83.000 48.800 85.000 49.100 ;
        RECT 6.200 48.100 6.600 48.200 ;
        RECT 12.600 48.100 13.000 48.200 ;
        RECT 6.200 47.800 13.000 48.100 ;
        RECT 14.200 48.100 14.600 48.200 ;
        RECT 17.400 48.100 17.800 48.200 ;
        RECT 14.200 47.800 17.800 48.100 ;
        RECT 18.200 48.100 18.600 48.200 ;
        RECT 20.600 48.100 21.000 48.200 ;
        RECT 18.200 47.800 21.000 48.100 ;
        RECT 23.000 48.100 23.400 48.200 ;
        RECT 29.400 48.100 29.800 48.200 ;
        RECT 23.000 47.800 29.800 48.100 ;
        RECT 52.600 48.100 53.000 48.200 ;
        RECT 57.400 48.100 57.800 48.200 ;
        RECT 52.600 47.800 57.800 48.100 ;
        RECT 78.200 48.100 78.600 48.200 ;
        RECT 79.800 48.100 80.200 48.200 ;
        RECT 78.200 47.800 80.200 48.100 ;
        RECT 11.000 47.100 11.400 47.200 ;
        RECT 11.000 46.800 12.100 47.100 ;
        RECT 11.800 46.200 12.100 46.800 ;
        RECT 15.000 46.800 15.400 47.200 ;
        RECT 22.200 47.100 22.600 47.200 ;
        RECT 15.800 46.800 22.600 47.100 ;
        RECT 23.800 47.100 24.200 47.200 ;
        RECT 28.600 47.100 29.000 47.200 ;
        RECT 23.800 46.800 29.000 47.100 ;
        RECT 30.200 47.100 30.600 47.200 ;
        RECT 31.000 47.100 31.400 47.200 ;
        RECT 30.200 46.800 31.400 47.100 ;
        RECT 35.000 47.100 35.400 47.200 ;
        RECT 35.800 47.100 36.200 47.200 ;
        RECT 35.000 46.800 36.200 47.100 ;
        RECT 42.200 47.100 42.600 47.200 ;
        RECT 52.600 47.100 53.000 47.200 ;
        RECT 42.200 46.800 53.000 47.100 ;
        RECT 84.600 47.100 85.000 47.200 ;
        RECT 86.200 47.100 86.600 47.200 ;
        RECT 84.600 46.800 86.600 47.100 ;
        RECT 15.000 46.200 15.300 46.800 ;
        RECT 15.800 46.200 16.100 46.800 ;
        RECT 3.000 46.100 3.400 46.200 ;
        RECT 7.000 46.100 7.400 46.200 ;
        RECT 3.000 45.800 7.400 46.100 ;
        RECT 10.200 46.100 10.600 46.200 ;
        RECT 11.000 46.100 11.400 46.200 ;
        RECT 10.200 45.800 11.400 46.100 ;
        RECT 11.800 45.800 12.200 46.200 ;
        RECT 15.000 45.800 15.400 46.200 ;
        RECT 15.800 45.800 16.200 46.200 ;
        RECT 16.600 46.100 17.000 46.200 ;
        RECT 20.600 46.100 21.000 46.200 ;
        RECT 16.600 45.800 21.000 46.100 ;
        RECT 27.800 45.800 28.200 46.200 ;
        RECT 31.800 46.100 32.200 46.200 ;
        RECT 30.200 45.800 32.200 46.100 ;
        RECT 39.000 45.800 39.400 46.200 ;
        RECT 45.400 46.100 45.800 46.200 ;
        RECT 47.000 46.100 47.400 46.200 ;
        RECT 45.400 45.800 47.400 46.100 ;
        RECT 50.200 46.100 50.600 46.200 ;
        RECT 63.800 46.100 64.200 46.200 ;
        RECT 67.000 46.100 67.400 46.200 ;
        RECT 50.200 45.800 67.400 46.100 ;
        RECT 71.800 46.100 72.200 46.200 ;
        RECT 74.200 46.100 74.600 46.200 ;
        RECT 71.800 45.800 74.600 46.100 ;
        RECT 79.000 46.100 79.400 46.200 ;
        RECT 81.400 46.100 81.800 46.200 ;
        RECT 79.000 45.800 81.800 46.100 ;
        RECT 6.200 45.100 6.600 45.200 ;
        RECT 7.000 45.100 7.400 45.200 ;
        RECT 6.200 44.800 7.400 45.100 ;
        RECT 11.800 45.100 12.200 45.200 ;
        RECT 19.800 45.100 20.200 45.200 ;
        RECT 11.800 44.800 20.200 45.100 ;
        RECT 26.200 45.100 26.600 45.200 ;
        RECT 27.800 45.100 28.100 45.800 ;
        RECT 26.200 44.800 28.100 45.100 ;
        RECT 30.200 45.200 30.500 45.800 ;
        RECT 30.200 44.800 30.600 45.200 ;
        RECT 31.000 45.100 31.400 45.200 ;
        RECT 32.600 45.100 33.000 45.200 ;
        RECT 39.000 45.100 39.300 45.800 ;
        RECT 31.000 44.800 39.300 45.100 ;
        RECT 54.200 45.100 54.600 45.200 ;
        RECT 72.600 45.100 73.000 45.200 ;
        RECT 77.400 45.100 77.800 45.200 ;
        RECT 54.200 44.800 77.800 45.100 ;
        RECT 75.000 44.100 75.400 44.200 ;
        RECT 78.200 44.100 78.600 44.200 ;
        RECT 75.000 43.800 78.600 44.100 ;
        RECT 9.400 43.100 9.800 43.200 ;
        RECT 10.200 43.100 10.600 43.200 ;
        RECT 42.200 43.100 42.600 43.200 ;
        RECT 77.400 43.100 77.800 43.200 ;
        RECT 79.000 43.100 79.400 43.200 ;
        RECT 9.400 42.800 79.400 43.100 ;
        RECT 30.200 42.100 30.600 42.200 ;
        RECT 31.000 42.100 31.400 42.200 ;
        RECT 30.200 41.800 31.400 42.100 ;
        RECT 59.800 42.100 60.200 42.200 ;
        RECT 74.200 42.100 74.600 42.200 ;
        RECT 75.800 42.100 76.200 42.200 ;
        RECT 59.800 41.800 76.200 42.100 ;
        RECT 62.200 41.100 62.600 41.200 ;
        RECT 71.800 41.100 72.200 41.200 ;
        RECT 62.200 40.800 72.200 41.100 ;
        RECT 47.800 40.100 48.200 40.200 ;
        RECT 67.800 40.100 68.200 40.200 ;
        RECT 47.800 39.800 68.200 40.100 ;
        RECT 82.200 40.100 82.600 40.200 ;
        RECT 83.800 40.100 84.200 40.200 ;
        RECT 82.200 39.800 84.200 40.100 ;
        RECT 21.400 39.100 21.800 39.200 ;
        RECT 25.400 39.100 25.800 39.200 ;
        RECT 55.800 39.100 56.200 39.200 ;
        RECT 56.600 39.100 57.000 39.200 ;
        RECT 21.400 38.800 57.000 39.100 ;
        RECT 18.200 38.100 18.600 38.200 ;
        RECT 43.000 38.100 43.400 38.200 ;
        RECT 18.200 37.800 43.400 38.100 ;
        RECT 55.800 37.800 56.200 38.200 ;
        RECT 56.600 38.100 57.000 38.200 ;
        RECT 69.400 38.100 69.800 38.200 ;
        RECT 81.400 38.100 81.800 38.200 ;
        RECT 84.600 38.100 85.000 38.200 ;
        RECT 56.600 37.800 85.000 38.100 ;
        RECT 3.800 37.100 4.200 37.200 ;
        RECT 12.600 37.100 13.000 37.200 ;
        RECT 3.800 36.800 13.000 37.100 ;
        RECT 25.400 37.100 25.800 37.200 ;
        RECT 27.000 37.100 27.400 37.200 ;
        RECT 25.400 36.800 27.400 37.100 ;
        RECT 55.800 37.100 56.100 37.800 ;
        RECT 67.000 37.100 67.400 37.200 ;
        RECT 55.800 36.800 67.400 37.100 ;
        RECT 74.200 36.800 74.600 37.200 ;
        RECT 80.600 37.100 81.000 37.200 ;
        RECT 80.600 36.800 82.500 37.100 ;
        RECT 6.200 36.100 6.600 36.200 ;
        RECT 7.000 36.100 7.400 36.200 ;
        RECT 6.200 35.800 7.400 36.100 ;
        RECT 7.800 36.100 8.200 36.200 ;
        RECT 11.800 36.100 12.200 36.200 ;
        RECT 7.800 35.800 12.200 36.100 ;
        RECT 20.600 36.100 21.000 36.200 ;
        RECT 23.800 36.100 24.200 36.200 ;
        RECT 20.600 35.800 24.200 36.100 ;
        RECT 28.600 36.100 29.000 36.200 ;
        RECT 40.600 36.100 41.000 36.200 ;
        RECT 44.600 36.100 45.000 36.200 ;
        RECT 28.600 35.800 31.300 36.100 ;
        RECT 40.600 35.800 45.000 36.100 ;
        RECT 57.400 36.100 57.800 36.200 ;
        RECT 58.200 36.100 58.600 36.200 ;
        RECT 57.400 35.800 58.600 36.100 ;
        RECT 68.600 36.100 69.000 36.200 ;
        RECT 74.200 36.100 74.500 36.800 ;
        RECT 68.600 35.800 74.500 36.100 ;
        RECT 82.200 36.200 82.500 36.800 ;
        RECT 82.200 35.800 82.600 36.200 ;
        RECT 31.000 35.200 31.300 35.800 ;
        RECT 9.400 35.100 9.800 35.200 ;
        RECT 15.800 35.100 16.200 35.200 ;
        RECT 21.400 35.100 21.800 35.200 ;
        RECT 9.400 34.800 21.800 35.100 ;
        RECT 31.000 34.800 31.400 35.200 ;
        RECT 48.600 35.100 49.000 35.200 ;
        RECT 51.000 35.100 51.400 35.200 ;
        RECT 48.600 34.800 51.400 35.100 ;
        RECT 53.400 35.100 53.800 35.200 ;
        RECT 54.200 35.100 54.600 35.200 ;
        RECT 53.400 34.800 54.600 35.100 ;
        RECT 55.000 35.100 55.400 35.200 ;
        RECT 55.800 35.100 56.200 35.200 ;
        RECT 55.000 34.800 56.200 35.100 ;
        RECT 58.200 35.100 58.600 35.200 ;
        RECT 59.000 35.100 59.400 35.200 ;
        RECT 58.200 34.800 59.400 35.100 ;
        RECT 60.600 35.100 61.000 35.200 ;
        RECT 65.400 35.100 65.800 35.200 ;
        RECT 60.600 34.800 65.800 35.100 ;
        RECT 67.800 35.100 68.200 35.200 ;
        RECT 74.200 35.100 74.600 35.200 ;
        RECT 75.800 35.100 76.200 35.200 ;
        RECT 67.800 34.800 73.700 35.100 ;
        RECT 74.200 34.800 76.200 35.100 ;
        RECT 82.200 35.100 82.600 35.200 ;
        RECT 85.400 35.100 85.800 35.200 ;
        RECT 82.200 34.800 85.800 35.100 ;
        RECT 6.200 34.100 6.600 34.200 ;
        RECT 9.400 34.100 9.700 34.800 ;
        RECT 6.200 33.800 9.700 34.100 ;
        RECT 11.000 34.100 11.400 34.200 ;
        RECT 17.400 34.100 17.800 34.200 ;
        RECT 11.000 33.800 17.800 34.100 ;
        RECT 19.000 34.100 19.400 34.200 ;
        RECT 51.000 34.100 51.400 34.200 ;
        RECT 19.000 33.800 51.400 34.100 ;
        RECT 58.200 34.100 58.600 34.200 ;
        RECT 67.800 34.100 68.200 34.200 ;
        RECT 68.600 34.100 69.000 34.200 ;
        RECT 58.200 33.800 69.000 34.100 ;
        RECT 69.400 34.100 69.800 34.200 ;
        RECT 71.800 34.100 72.200 34.200 ;
        RECT 69.400 33.800 72.200 34.100 ;
        RECT 73.400 34.100 73.700 34.800 ;
        RECT 79.000 34.100 79.400 34.200 ;
        RECT 73.400 33.800 79.400 34.100 ;
        RECT 79.800 34.100 80.200 34.200 ;
        RECT 84.600 34.100 85.000 34.200 ;
        RECT 79.800 33.800 85.000 34.100 ;
        RECT 8.600 33.100 9.000 33.200 ;
        RECT 11.800 33.100 12.200 33.200 ;
        RECT 8.600 32.800 12.200 33.100 ;
        RECT 14.200 32.800 14.600 33.200 ;
        RECT 28.600 33.100 29.000 33.200 ;
        RECT 26.200 32.800 29.000 33.100 ;
        RECT 34.200 33.100 34.600 33.200 ;
        RECT 35.000 33.100 35.400 33.200 ;
        RECT 36.600 33.100 37.000 33.200 ;
        RECT 34.200 32.800 37.000 33.100 ;
        RECT 38.200 33.100 38.600 33.200 ;
        RECT 40.600 33.100 41.000 33.200 ;
        RECT 51.800 33.100 52.200 33.200 ;
        RECT 38.200 32.800 41.000 33.100 ;
        RECT 45.400 32.800 52.200 33.100 ;
        RECT 54.200 33.100 54.600 33.200 ;
        RECT 59.800 33.100 60.200 33.200 ;
        RECT 54.200 32.800 60.200 33.100 ;
        RECT 67.000 33.100 67.400 33.200 ;
        RECT 67.800 33.100 68.200 33.200 ;
        RECT 67.000 32.800 68.200 33.100 ;
        RECT 14.200 32.100 14.500 32.800 ;
        RECT 26.200 32.200 26.500 32.800 ;
        RECT 45.400 32.200 45.700 32.800 ;
        RECT 24.600 32.100 25.000 32.200 ;
        RECT 14.200 31.800 25.000 32.100 ;
        RECT 26.200 32.100 26.600 32.200 ;
        RECT 35.800 32.100 36.200 32.200 ;
        RECT 26.200 31.800 36.200 32.100 ;
        RECT 38.200 32.100 38.600 32.200 ;
        RECT 39.800 32.100 40.200 32.200 ;
        RECT 38.200 31.800 40.200 32.100 ;
        RECT 44.600 32.100 45.000 32.200 ;
        RECT 45.400 32.100 45.800 32.200 ;
        RECT 44.600 31.800 45.800 32.100 ;
        RECT 46.200 32.100 46.600 32.200 ;
        RECT 47.000 32.100 47.400 32.200 ;
        RECT 59.000 32.100 59.400 32.200 ;
        RECT 64.600 32.100 65.000 32.200 ;
        RECT 46.200 31.800 47.400 32.100 ;
        RECT 58.200 31.800 65.000 32.100 ;
        RECT 77.400 31.800 77.800 32.200 ;
        RECT 77.400 31.200 77.700 31.800 ;
        RECT 6.200 31.100 6.600 31.200 ;
        RECT 8.600 31.100 9.000 31.200 ;
        RECT 20.600 31.100 21.000 31.200 ;
        RECT 6.200 30.800 21.000 31.100 ;
        RECT 50.200 31.100 50.600 31.200 ;
        RECT 59.800 31.100 60.200 31.200 ;
        RECT 50.200 30.800 60.200 31.100 ;
        RECT 77.400 30.800 77.800 31.200 ;
        RECT 36.600 30.100 37.000 30.200 ;
        RECT 49.400 30.100 49.800 30.200 ;
        RECT 36.600 29.800 49.800 30.100 ;
        RECT 74.200 30.100 74.600 30.200 ;
        RECT 77.400 30.100 77.800 30.200 ;
        RECT 74.200 29.800 77.800 30.100 ;
        RECT 6.200 29.100 6.600 29.200 ;
        RECT 11.800 29.100 12.200 29.200 ;
        RECT 6.200 28.800 12.200 29.100 ;
        RECT 18.200 29.100 18.600 29.200 ;
        RECT 22.200 29.100 22.600 29.200 ;
        RECT 18.200 28.800 22.600 29.100 ;
        RECT 31.800 29.100 32.200 29.200 ;
        RECT 33.400 29.100 33.800 29.200 ;
        RECT 44.600 29.100 45.000 29.200 ;
        RECT 31.800 28.800 33.800 29.100 ;
        RECT 35.000 28.800 45.000 29.100 ;
        RECT 49.400 29.100 49.800 29.200 ;
        RECT 51.800 29.100 52.200 29.200 ;
        RECT 72.600 29.100 73.000 29.200 ;
        RECT 49.400 28.800 52.200 29.100 ;
        RECT 52.600 28.800 73.000 29.100 ;
        RECT 35.000 28.200 35.300 28.800 ;
        RECT 7.800 28.100 8.200 28.200 ;
        RECT 14.200 28.100 14.600 28.200 ;
        RECT 7.800 27.800 14.600 28.100 ;
        RECT 16.600 28.100 17.000 28.200 ;
        RECT 19.800 28.100 20.200 28.200 ;
        RECT 16.600 27.800 20.200 28.100 ;
        RECT 20.600 28.100 21.000 28.200 ;
        RECT 21.400 28.100 21.800 28.200 ;
        RECT 20.600 27.800 21.800 28.100 ;
        RECT 35.000 27.800 35.400 28.200 ;
        RECT 35.800 28.100 36.200 28.200 ;
        RECT 43.000 28.100 43.400 28.200 ;
        RECT 35.800 27.800 43.400 28.100 ;
        RECT 50.200 28.100 50.600 28.200 ;
        RECT 52.600 28.100 52.900 28.800 ;
        RECT 50.200 27.800 52.900 28.100 ;
        RECT 63.800 28.100 64.200 28.200 ;
        RECT 68.600 28.100 69.000 28.200 ;
        RECT 63.800 27.800 69.000 28.100 ;
        RECT 69.400 28.100 69.800 28.200 ;
        RECT 73.400 28.100 73.800 28.200 ;
        RECT 81.400 28.100 81.800 28.200 ;
        RECT 69.400 27.800 81.800 28.100 ;
        RECT 37.400 27.100 37.800 27.200 ;
        RECT 39.000 27.100 39.400 27.200 ;
        RECT 37.400 26.800 39.400 27.100 ;
        RECT 53.400 27.100 53.800 27.200 ;
        RECT 55.800 27.100 56.200 27.200 ;
        RECT 53.400 26.800 56.200 27.100 ;
        RECT 58.200 27.100 58.600 27.200 ;
        RECT 64.600 27.100 65.000 27.200 ;
        RECT 58.200 26.800 65.000 27.100 ;
        RECT 67.800 27.100 68.200 27.200 ;
        RECT 72.600 27.100 73.000 27.200 ;
        RECT 67.800 26.800 73.000 27.100 ;
        RECT 75.800 27.100 76.200 27.200 ;
        RECT 76.600 27.100 77.000 27.200 ;
        RECT 75.800 26.800 77.000 27.100 ;
        RECT 10.200 26.100 10.600 26.200 ;
        RECT 19.800 26.100 20.200 26.200 ;
        RECT 10.200 25.800 20.200 26.100 ;
        RECT 23.000 26.100 23.400 26.200 ;
        RECT 32.600 26.100 33.000 26.200 ;
        RECT 39.800 26.100 40.200 26.200 ;
        RECT 23.000 25.800 40.200 26.100 ;
        RECT 47.800 26.100 48.200 26.200 ;
        RECT 54.200 26.100 54.600 26.200 ;
        RECT 55.000 26.100 55.400 26.200 ;
        RECT 47.800 25.800 50.500 26.100 ;
        RECT 54.200 25.800 55.400 26.100 ;
        RECT 63.800 26.100 64.200 26.200 ;
        RECT 66.200 26.100 66.600 26.200 ;
        RECT 71.000 26.100 71.400 26.200 ;
        RECT 84.600 26.100 85.000 26.200 ;
        RECT 63.800 25.800 85.000 26.100 ;
        RECT 7.000 25.100 7.400 25.200 ;
        RECT 9.400 25.100 9.800 25.200 ;
        RECT 7.000 24.800 9.800 25.100 ;
        RECT 15.000 25.100 15.400 25.200 ;
        RECT 45.400 25.100 45.800 25.200 ;
        RECT 49.400 25.100 49.800 25.200 ;
        RECT 15.000 24.800 49.800 25.100 ;
        RECT 50.200 25.100 50.500 25.800 ;
        RECT 61.400 25.100 61.800 25.200 ;
        RECT 82.200 25.100 82.600 25.200 ;
        RECT 50.200 24.800 67.300 25.100 ;
        RECT 67.000 24.200 67.300 24.800 ;
        RECT 79.800 24.800 82.600 25.100 ;
        RECT 79.800 24.200 80.100 24.800 ;
        RECT 13.400 24.100 13.800 24.200 ;
        RECT 41.400 24.100 41.800 24.200 ;
        RECT 13.400 23.800 41.800 24.100 ;
        RECT 47.800 24.100 48.200 24.200 ;
        RECT 51.000 24.100 51.400 24.200 ;
        RECT 47.800 23.800 51.400 24.100 ;
        RECT 67.000 23.800 67.400 24.200 ;
        RECT 79.800 23.800 80.200 24.200 ;
        RECT 14.200 23.100 14.600 23.200 ;
        RECT 31.000 23.100 31.400 23.200 ;
        RECT 14.200 22.800 31.400 23.100 ;
        RECT 15.000 22.100 15.400 22.200 ;
        RECT 33.400 22.100 33.800 22.200 ;
        RECT 15.000 21.800 33.800 22.100 ;
        RECT 51.000 22.100 51.400 22.200 ;
        RECT 80.600 22.100 81.000 22.200 ;
        RECT 85.400 22.100 85.800 22.200 ;
        RECT 51.000 21.800 85.800 22.100 ;
        RECT 67.000 21.100 67.400 21.200 ;
        RECT 69.400 21.100 69.800 21.200 ;
        RECT 83.000 21.100 83.400 21.200 ;
        RECT 67.000 20.800 83.400 21.100 ;
        RECT 44.600 20.100 45.000 20.200 ;
        RECT 65.400 20.100 65.800 20.200 ;
        RECT 80.600 20.100 81.000 20.200 ;
        RECT 44.600 19.800 81.000 20.100 ;
        RECT 5.400 19.100 5.800 19.200 ;
        RECT 9.400 19.100 9.800 19.200 ;
        RECT 5.400 18.800 9.800 19.100 ;
        RECT 14.200 19.100 14.600 19.200 ;
        RECT 18.200 19.100 18.600 19.200 ;
        RECT 14.200 18.800 18.600 19.100 ;
        RECT 55.800 19.100 56.200 19.200 ;
        RECT 71.800 19.100 72.200 19.200 ;
        RECT 55.800 18.800 72.200 19.100 ;
        RECT 3.800 18.100 4.200 18.200 ;
        RECT 6.200 18.100 6.600 18.200 ;
        RECT 11.000 18.100 11.400 18.200 ;
        RECT 13.400 18.100 13.800 18.200 ;
        RECT 3.800 17.800 13.800 18.100 ;
        RECT 18.200 18.100 18.600 18.200 ;
        RECT 20.600 18.100 21.000 18.200 ;
        RECT 18.200 17.800 21.000 18.100 ;
        RECT 25.400 18.100 25.800 18.200 ;
        RECT 54.200 18.100 54.600 18.200 ;
        RECT 25.400 17.800 54.600 18.100 ;
        RECT 57.400 17.800 57.800 18.200 ;
        RECT 9.400 17.100 9.800 17.200 ;
        RECT 19.000 17.100 19.400 17.200 ;
        RECT 9.400 16.800 19.400 17.100 ;
        RECT 22.200 16.800 22.600 17.200 ;
        RECT 32.600 16.800 33.000 17.200 ;
        RECT 45.400 17.100 45.800 17.200 ;
        RECT 57.400 17.100 57.700 17.800 ;
        RECT 45.400 16.800 57.700 17.100 ;
        RECT 3.800 16.100 4.200 16.200 ;
        RECT 22.200 16.100 22.500 16.800 ;
        RECT 3.800 15.800 22.500 16.100 ;
        RECT 23.000 16.100 23.400 16.200 ;
        RECT 32.600 16.100 32.900 16.800 ;
        RECT 23.000 15.800 32.900 16.100 ;
        RECT 36.600 16.100 37.000 16.200 ;
        RECT 38.200 16.100 38.600 16.200 ;
        RECT 36.600 15.800 38.600 16.100 ;
        RECT 44.600 16.100 45.000 16.200 ;
        RECT 46.200 16.100 46.600 16.200 ;
        RECT 44.600 15.800 46.600 16.100 ;
        RECT 47.800 16.100 48.200 16.200 ;
        RECT 52.600 16.100 53.000 16.200 ;
        RECT 47.800 15.800 53.000 16.100 ;
        RECT 53.400 16.100 53.800 16.200 ;
        RECT 55.000 16.100 55.400 16.200 ;
        RECT 68.600 16.100 69.000 16.200 ;
        RECT 53.400 15.800 55.400 16.100 ;
        RECT 66.200 15.800 69.000 16.100 ;
        RECT 80.600 16.100 81.000 16.200 ;
        RECT 83.000 16.100 83.400 16.200 ;
        RECT 80.600 15.800 83.400 16.100 ;
        RECT 66.200 15.200 66.500 15.800 ;
        RECT 5.400 15.100 5.800 15.200 ;
        RECT 7.000 15.100 7.400 15.200 ;
        RECT 5.400 14.800 7.400 15.100 ;
        RECT 15.800 15.100 16.200 15.200 ;
        RECT 16.600 15.100 17.000 15.200 ;
        RECT 15.800 14.800 17.000 15.100 ;
        RECT 20.600 15.100 21.000 15.200 ;
        RECT 23.800 15.100 24.200 15.200 ;
        RECT 20.600 14.800 24.200 15.100 ;
        RECT 31.800 15.100 32.200 15.200 ;
        RECT 32.600 15.100 33.000 15.200 ;
        RECT 41.400 15.100 41.800 15.200 ;
        RECT 49.400 15.100 49.800 15.200 ;
        RECT 56.600 15.100 57.000 15.200 ;
        RECT 31.800 14.800 57.000 15.100 ;
        RECT 58.200 15.100 58.600 15.200 ;
        RECT 62.200 15.100 62.600 15.200 ;
        RECT 58.200 14.800 62.600 15.100 ;
        RECT 66.200 14.800 66.600 15.200 ;
        RECT 71.000 15.100 71.400 15.200 ;
        RECT 77.400 15.100 77.800 15.200 ;
        RECT 80.600 15.100 81.000 15.200 ;
        RECT 71.000 14.800 81.000 15.100 ;
        RECT 83.000 15.100 83.400 15.200 ;
        RECT 84.600 15.100 85.000 15.200 ;
        RECT 83.000 14.800 85.000 15.100 ;
        RECT 7.000 14.100 7.400 14.200 ;
        RECT 12.600 14.100 13.000 14.200 ;
        RECT 7.000 13.800 13.000 14.100 ;
        RECT 31.000 13.800 31.400 14.200 ;
        RECT 35.800 13.800 36.200 14.200 ;
        RECT 36.600 14.100 37.000 14.200 ;
        RECT 39.000 14.100 39.400 14.200 ;
        RECT 45.400 14.100 45.800 14.200 ;
        RECT 36.600 13.800 39.400 14.100 ;
        RECT 43.800 13.800 45.800 14.100 ;
        RECT 52.600 14.100 53.000 14.200 ;
        RECT 53.400 14.100 53.800 14.200 ;
        RECT 52.600 13.800 53.800 14.100 ;
        RECT 54.200 14.100 54.600 14.200 ;
        RECT 67.000 14.100 67.400 14.200 ;
        RECT 54.200 13.800 67.400 14.100 ;
        RECT 77.400 14.100 77.800 14.200 ;
        RECT 79.800 14.100 80.200 14.200 ;
        RECT 77.400 13.800 80.200 14.100 ;
        RECT 82.200 14.100 82.600 14.200 ;
        RECT 83.000 14.100 83.400 14.200 ;
        RECT 82.200 13.800 83.400 14.100 ;
        RECT 18.200 13.100 18.600 13.200 ;
        RECT 19.800 13.100 20.200 13.200 ;
        RECT 18.200 12.800 20.200 13.100 ;
        RECT 31.000 13.100 31.300 13.800 ;
        RECT 35.800 13.100 36.100 13.800 ;
        RECT 31.000 12.800 36.100 13.100 ;
        RECT 43.800 13.200 44.100 13.800 ;
        RECT 43.800 12.800 44.200 13.200 ;
        RECT 47.800 13.100 48.200 13.200 ;
        RECT 49.400 13.100 49.800 13.200 ;
        RECT 47.800 12.800 49.800 13.100 ;
        RECT 53.400 13.100 53.700 13.800 ;
        RECT 69.400 13.100 69.800 13.200 ;
        RECT 53.400 12.800 69.800 13.100 ;
        RECT 71.800 13.100 72.200 13.200 ;
        RECT 75.000 13.100 75.400 13.200 ;
        RECT 71.800 12.800 75.400 13.100 ;
        RECT 83.800 13.100 84.200 13.200 ;
        RECT 84.600 13.100 85.000 13.200 ;
        RECT 83.800 12.800 85.000 13.100 ;
        RECT 31.800 12.100 32.200 12.200 ;
        RECT 38.200 12.100 38.600 12.200 ;
        RECT 48.600 12.100 49.000 12.200 ;
        RECT 31.800 11.800 49.000 12.100 ;
        RECT 55.800 12.100 56.200 12.200 ;
        RECT 58.200 12.100 58.600 12.200 ;
        RECT 59.800 12.100 60.200 12.200 ;
        RECT 64.600 12.100 65.000 12.200 ;
        RECT 67.000 12.100 67.400 12.200 ;
        RECT 71.000 12.100 71.400 12.200 ;
        RECT 74.200 12.100 74.600 12.200 ;
        RECT 76.600 12.100 77.000 12.200 ;
        RECT 55.800 11.800 65.000 12.100 ;
        RECT 66.200 11.800 71.400 12.100 ;
        RECT 73.400 11.800 77.000 12.100 ;
        RECT 23.800 11.100 24.200 11.200 ;
        RECT 39.800 11.100 40.200 11.200 ;
        RECT 23.800 10.800 40.200 11.100 ;
        RECT 41.400 11.100 41.800 11.200 ;
        RECT 51.000 11.100 51.400 11.200 ;
        RECT 41.400 10.800 51.400 11.100 ;
        RECT 52.600 11.100 53.000 11.200 ;
        RECT 55.000 11.100 55.400 11.200 ;
        RECT 59.000 11.100 59.400 11.200 ;
        RECT 52.600 10.800 59.400 11.100 ;
        RECT 75.800 11.100 76.200 11.200 ;
        RECT 83.800 11.100 84.200 11.200 ;
        RECT 75.800 10.800 84.200 11.100 ;
        RECT 13.400 10.100 13.800 10.200 ;
        RECT 16.600 10.100 17.000 10.200 ;
        RECT 13.400 9.800 17.000 10.100 ;
        RECT 34.200 10.100 34.600 10.200 ;
        RECT 37.400 10.100 37.800 10.200 ;
        RECT 34.200 9.800 37.800 10.100 ;
        RECT 44.600 10.100 45.000 10.200 ;
        RECT 45.400 10.100 45.800 10.200 ;
        RECT 44.600 9.800 45.800 10.100 ;
        RECT 73.400 10.100 73.800 10.200 ;
        RECT 77.400 10.100 77.800 10.200 ;
        RECT 79.000 10.100 79.400 10.200 ;
        RECT 73.400 9.800 79.400 10.100 ;
        RECT 7.800 9.100 8.200 9.200 ;
        RECT 18.200 9.100 18.600 9.200 ;
        RECT 7.800 8.800 18.600 9.100 ;
        RECT 41.400 8.800 41.800 9.200 ;
        RECT 43.800 9.100 44.200 9.200 ;
        RECT 47.000 9.100 47.400 9.200 ;
        RECT 51.800 9.100 52.200 9.200 ;
        RECT 63.000 9.100 63.400 9.200 ;
        RECT 43.800 8.800 63.400 9.100 ;
        RECT 67.800 9.100 68.200 9.200 ;
        RECT 78.200 9.100 78.600 9.200 ;
        RECT 67.800 8.800 78.600 9.100 ;
        RECT 3.000 7.800 3.400 8.200 ;
        RECT 41.400 8.100 41.700 8.800 ;
        RECT 46.200 8.100 46.600 8.200 ;
        RECT 41.400 7.800 46.600 8.100 ;
        RECT 51.000 8.100 51.400 8.200 ;
        RECT 54.200 8.100 54.600 8.200 ;
        RECT 60.600 8.100 61.000 8.200 ;
        RECT 51.000 7.800 61.000 8.100 ;
        RECT 63.000 8.100 63.400 8.200 ;
        RECT 66.200 8.100 66.600 8.200 ;
        RECT 63.000 7.800 66.600 8.100 ;
        RECT 3.000 7.100 3.300 7.800 ;
        RECT 15.000 7.100 15.400 7.200 ;
        RECT 3.000 6.800 15.400 7.100 ;
        RECT 37.400 7.100 37.800 7.200 ;
        RECT 42.200 7.100 42.600 7.200 ;
        RECT 37.400 6.800 42.600 7.100 ;
        RECT 47.800 7.100 48.200 7.200 ;
        RECT 61.400 7.100 61.800 7.200 ;
        RECT 63.000 7.100 63.400 7.200 ;
        RECT 47.800 6.800 53.700 7.100 ;
        RECT 61.400 6.800 63.400 7.100 ;
        RECT 3.000 6.100 3.400 6.200 ;
        RECT 10.200 6.100 10.600 6.200 ;
        RECT 3.000 5.800 10.600 6.100 ;
        RECT 39.800 6.100 40.200 6.200 ;
        RECT 41.400 6.100 41.800 6.200 ;
        RECT 39.800 5.800 41.800 6.100 ;
        RECT 42.200 5.800 42.600 6.200 ;
        RECT 50.200 6.100 50.600 6.200 ;
        RECT 52.600 6.100 53.000 6.200 ;
        RECT 50.200 5.800 53.000 6.100 ;
        RECT 53.400 6.100 53.700 6.800 ;
        RECT 74.200 6.100 74.600 6.200 ;
        RECT 53.400 5.800 74.600 6.100 ;
        RECT 79.800 6.100 80.200 6.200 ;
        RECT 81.400 6.100 81.800 6.200 ;
        RECT 79.800 5.800 81.800 6.100 ;
        RECT 42.200 5.200 42.500 5.800 ;
        RECT 42.200 4.800 42.600 5.200 ;
        RECT 64.600 5.100 65.000 5.200 ;
        RECT 67.000 5.100 67.400 5.200 ;
        RECT 64.600 4.800 67.400 5.100 ;
      LAYER via3 ;
        RECT 54.200 64.800 54.600 65.200 ;
        RECT 84.600 58.800 85.000 59.200 ;
        RECT 83.000 57.800 83.400 58.200 ;
        RECT 11.000 56.800 11.400 57.200 ;
        RECT 53.400 55.800 53.800 56.200 ;
        RECT 75.000 51.800 75.400 52.200 ;
        RECT 35.800 50.800 36.200 51.200 ;
        RECT 57.400 50.800 57.800 51.200 ;
        RECT 31.000 46.800 31.400 47.200 ;
        RECT 11.000 45.800 11.400 46.200 ;
        RECT 32.600 44.800 33.000 45.200 ;
        RECT 42.200 42.800 42.600 43.200 ;
        RECT 31.000 41.800 31.400 42.200 ;
        RECT 67.800 39.800 68.200 40.200 ;
        RECT 55.800 38.800 56.200 39.200 ;
        RECT 58.200 35.800 58.600 36.200 ;
        RECT 51.000 34.800 51.400 35.200 ;
        RECT 54.200 34.800 54.600 35.200 ;
        RECT 55.800 34.800 56.200 35.200 ;
        RECT 68.600 33.800 69.000 34.200 ;
        RECT 35.000 32.800 35.400 33.200 ;
        RECT 24.600 31.800 25.000 32.200 ;
        RECT 21.400 27.800 21.800 28.200 ;
        RECT 76.600 26.800 77.000 27.200 ;
        RECT 49.400 24.800 49.800 25.200 ;
        RECT 80.600 21.800 81.000 22.200 ;
        RECT 83.000 20.800 83.400 21.200 ;
        RECT 6.200 17.800 6.600 18.200 ;
        RECT 32.600 14.800 33.000 15.200 ;
        RECT 83.000 13.800 83.400 14.200 ;
        RECT 84.600 12.800 85.000 13.200 ;
        RECT 45.400 9.800 45.800 10.200 ;
        RECT 54.200 7.800 54.600 8.200 ;
      LAYER metal4 ;
        RECT 80.600 65.800 81.000 66.200 ;
        RECT 54.200 64.800 54.600 65.200 ;
        RECT 11.000 56.800 11.400 57.200 ;
        RECT 6.200 47.800 6.600 48.200 ;
        RECT 6.200 45.200 6.500 47.800 ;
        RECT 11.000 46.200 11.300 56.800 ;
        RECT 53.400 55.800 53.800 56.200 ;
        RECT 35.800 50.800 36.200 51.200 ;
        RECT 15.000 47.100 15.400 47.200 ;
        RECT 15.800 47.100 16.200 47.200 ;
        RECT 15.000 46.800 16.200 47.100 ;
        RECT 23.000 47.100 23.400 47.200 ;
        RECT 23.800 47.100 24.200 47.200 ;
        RECT 23.000 46.800 24.200 47.100 ;
        RECT 31.000 46.800 31.400 47.200 ;
        RECT 35.000 46.800 35.400 47.200 ;
        RECT 11.000 45.800 11.400 46.200 ;
        RECT 6.200 44.800 6.600 45.200 ;
        RECT 31.000 42.200 31.300 46.800 ;
        RECT 32.600 44.800 33.000 45.200 ;
        RECT 31.000 41.800 31.400 42.200 ;
        RECT 21.400 38.800 21.800 39.200 ;
        RECT 6.200 35.800 6.600 36.200 ;
        RECT 6.200 18.200 6.500 35.800 ;
        RECT 21.400 28.200 21.700 38.800 ;
        RECT 24.600 32.100 25.000 32.200 ;
        RECT 25.400 32.100 25.800 32.200 ;
        RECT 24.600 31.800 25.800 32.100 ;
        RECT 21.400 27.800 21.800 28.200 ;
        RECT 6.200 17.800 6.600 18.200 ;
        RECT 32.600 15.200 32.900 44.800 ;
        RECT 35.000 33.200 35.300 46.800 ;
        RECT 35.000 32.800 35.400 33.200 ;
        RECT 35.800 28.200 36.100 50.800 ;
        RECT 52.600 47.800 53.000 48.200 ;
        RECT 42.200 42.800 42.600 43.200 ;
        RECT 35.800 27.800 36.200 28.200 ;
        RECT 15.800 15.100 16.200 15.200 ;
        RECT 16.600 15.100 17.000 15.200 ;
        RECT 15.800 14.800 17.000 15.100 ;
        RECT 32.600 14.800 33.000 15.200 ;
        RECT 36.600 14.800 37.000 15.200 ;
        RECT 36.600 14.200 36.900 14.800 ;
        RECT 36.600 13.800 37.000 14.200 ;
        RECT 42.200 5.200 42.500 42.800 ;
        RECT 51.000 35.100 51.400 35.200 ;
        RECT 51.800 35.100 52.200 35.200 ;
        RECT 51.000 34.800 52.200 35.100 ;
        RECT 44.600 31.800 45.000 32.200 ;
        RECT 46.200 32.100 46.600 32.200 ;
        RECT 47.000 32.100 47.400 32.200 ;
        RECT 46.200 31.800 47.400 32.100 ;
        RECT 44.600 10.100 44.900 31.800 ;
        RECT 49.400 26.800 49.800 27.200 ;
        RECT 49.400 25.200 49.700 26.800 ;
        RECT 49.400 24.800 49.800 25.200 ;
        RECT 52.600 14.200 52.900 47.800 ;
        RECT 53.400 27.200 53.700 55.800 ;
        RECT 54.200 45.200 54.500 64.800 ;
        RECT 75.000 52.100 75.400 52.200 ;
        RECT 74.200 51.800 75.400 52.100 ;
        RECT 57.400 50.800 57.800 51.200 ;
        RECT 54.200 44.800 54.600 45.200 ;
        RECT 55.800 38.800 56.200 39.200 ;
        RECT 55.800 35.200 56.100 38.800 ;
        RECT 57.400 36.100 57.700 50.800 ;
        RECT 67.800 39.800 68.200 40.200 ;
        RECT 58.200 36.100 58.600 36.200 ;
        RECT 57.400 35.800 58.600 36.100 ;
        RECT 54.200 34.800 54.600 35.200 ;
        RECT 55.800 34.800 56.200 35.200 ;
        RECT 58.200 35.100 58.600 35.200 ;
        RECT 59.000 35.100 59.400 35.200 ;
        RECT 58.200 34.800 59.400 35.100 ;
        RECT 54.200 34.200 54.500 34.800 ;
        RECT 54.200 33.800 54.600 34.200 ;
        RECT 57.400 34.100 57.800 34.200 ;
        RECT 58.200 34.100 58.600 34.200 ;
        RECT 57.400 33.800 58.600 34.100 ;
        RECT 67.800 27.200 68.100 39.800 ;
        RECT 68.600 35.800 69.000 36.200 ;
        RECT 68.600 34.200 68.900 35.800 ;
        RECT 68.600 33.800 69.000 34.200 ;
        RECT 74.200 30.200 74.500 51.800 ;
        RECT 77.400 30.800 77.800 31.200 ;
        RECT 74.200 29.800 74.600 30.200 ;
        RECT 53.400 26.800 53.800 27.200 ;
        RECT 67.800 26.800 68.200 27.200 ;
        RECT 75.800 27.100 76.200 27.200 ;
        RECT 76.600 27.100 77.000 27.200 ;
        RECT 75.800 26.800 77.000 27.100 ;
        RECT 54.200 25.800 54.600 26.200 ;
        RECT 52.600 13.800 53.000 14.200 ;
        RECT 45.400 10.100 45.800 10.200 ;
        RECT 44.600 9.800 45.800 10.100 ;
        RECT 54.200 8.200 54.500 25.800 ;
        RECT 77.400 14.200 77.700 30.800 ;
        RECT 80.600 22.200 80.900 65.800 ;
        RECT 84.600 58.800 85.000 59.200 ;
        RECT 83.000 57.800 83.400 58.200 ;
        RECT 80.600 21.800 81.000 22.200 ;
        RECT 83.000 21.200 83.300 57.800 ;
        RECT 83.000 20.800 83.400 21.200 ;
        RECT 83.000 14.200 83.300 20.800 ;
        RECT 77.400 13.800 77.800 14.200 ;
        RECT 83.000 13.800 83.400 14.200 ;
        RECT 84.600 13.200 84.900 58.800 ;
        RECT 84.600 12.800 85.000 13.200 ;
        RECT 54.200 7.800 54.600 8.200 ;
        RECT 42.200 4.800 42.600 5.200 ;
      LAYER via4 ;
        RECT 15.800 46.800 16.200 47.200 ;
        RECT 25.400 31.800 25.800 32.200 ;
        RECT 16.600 14.800 17.000 15.200 ;
        RECT 51.800 34.800 52.200 35.200 ;
        RECT 47.000 31.800 47.400 32.200 ;
        RECT 59.000 34.800 59.400 35.200 ;
      LAYER metal5 ;
        RECT 15.800 47.100 16.200 47.200 ;
        RECT 23.000 47.100 23.400 47.200 ;
        RECT 15.800 46.800 23.400 47.100 ;
        RECT 51.800 35.100 52.200 35.200 ;
        RECT 59.000 35.100 59.400 35.200 ;
        RECT 51.800 34.800 59.400 35.100 ;
        RECT 54.200 34.100 54.600 34.200 ;
        RECT 57.400 34.100 57.800 34.200 ;
        RECT 54.200 33.800 57.800 34.100 ;
        RECT 25.400 32.100 25.800 32.200 ;
        RECT 47.000 32.100 47.400 32.200 ;
        RECT 25.400 31.800 47.400 32.100 ;
        RECT 49.400 27.100 49.800 27.200 ;
        RECT 75.800 27.100 76.200 27.200 ;
        RECT 49.400 26.800 76.200 27.100 ;
        RECT 16.600 15.100 17.000 15.200 ;
        RECT 36.600 15.100 37.000 15.200 ;
        RECT 16.600 14.800 37.000 15.100 ;
  END
END ALU_8bit
END LIBRARY

