* NGSPICE file created from ALU_8bit.ext - technology: scmos

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

.subckt ALU_8bit vdd gnd A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] B[0] B[1] B[2] B[3]
+ B[4] B[5] B[6] B[7] ALU_Sel[0] ALU_Sel[1] ALU_Sel[2] ALU_Out[0] ALU_Out[1] ALU_Out[2]
+ ALU_Out[3] ALU_Out[4] ALU_Out[5] ALU_Out[6] ALU_Out[7] CarryOut
XAND2X2_5 AND2X2_5/A AND2X2_5/B gnd AND2X2_5/Y vdd AND2X2
XNAND2X1_21 INVX2_8/Y OAI21X1_9/Y gnd AOI22X1_2/A vdd NAND2X1
XNAND2X1_10 NOR2X1_26/A NOR2X1_26/B gnd OAI21X1_4/A vdd NAND2X1
XINVX2_12 INVX2_12/A gnd INVX2_12/Y vdd INVX2
XOAI21X1_19 INVX2_11/Y NAND2X1_9/Y OAI21X1_19/C gnd AND2X2_5/B vdd OAI21X1
XFILL_0_0_0 gnd vdd FILL
XINVX1_6 B[4] gnd INVX1_6/Y vdd INVX1
XXNOR2X1_6 XNOR2X1_6/A AND2X2_1/Y gnd XNOR2X1_6/Y vdd XNOR2X1
XNAND2X1_22 ALU_Sel[0] ALU_Sel[1] gnd OR2X2_1/A vdd NAND2X1
XAOI22X1_1 INVX2_13/A AND2X2_3/Y INVX2_8/Y INVX2_12/A gnd NAND3X1_2/C vdd AOI22X1
XAND2X2_6 AND2X2_6/A AND2X2_6/B gnd AND2X2_6/Y vdd AND2X2
XNAND2X1_11 B[3] INVX2_6/Y gnd AOI21X1_4/A vdd NAND2X1
XINVX2_13 INVX2_13/A gnd INVX2_13/Y vdd INVX2
XFILL_0_0_1 gnd vdd FILL
XAND2X2_7 AND2X2_7/A AND2X2_7/B gnd AND2X2_7/Y vdd AND2X2
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XAOI22X1_2 AOI22X1_2/A AOI22X1_2/B OAI21X1_6/Y INVX4_4/A gnd AOI22X1_2/Y vdd AOI22X1
XNAND2X1_23 INVX1_11/Y INVX2_1/Y gnd NOR2X1_16/B vdd NAND2X1
XNAND2X1_12 AND2X2_1/B AND2X2_1/A gnd NOR2X1_11/A vdd NAND2X1
XINVX1_8 B[1] gnd INVX1_8/Y vdd INVX1
XAOI22X1_3 INVX2_13/A INVX2_9/Y A[1] INVX4_3/A gnd AND2X2_4/B vdd AOI22X1
XAND2X2_8 AND2X2_8/A AND2X2_8/B gnd AND2X2_8/Y vdd AND2X2
XNAND2X1_24 ALU_Sel[1] INVX1_11/Y gnd NOR2X1_14/B vdd NAND2X1
XNAND2X1_13 A[4] B[4] gnd AND2X2_7/B vdd NAND2X1
XFILL_3_0_0 gnd vdd FILL
XINVX1_9 B[2] gnd INVX1_9/Y vdd INVX1
XNAND2X1_25 A[1] INVX1_8/Y gnd AOI21X1_9/A vdd NAND2X1
XAOI22X1_4 INVX2_13/A NOR2X1_9/Y A[0] INVX1_14/A gnd AOI22X1_4/Y vdd AOI22X1
XNAND2X1_14 INVX4_1/Y INVX1_6/Y gnd AND2X2_7/A vdd NAND2X1
XFILL_3_0_1 gnd vdd FILL
XAOI22X1_5 INVX2_13/A INVX1_12/A A[1] INVX1_14/A gnd AOI22X1_5/Y vdd AOI22X1
XNAND2X1_26 NOR2X1_26/B AOI21X1_6/Y gnd NAND3X1_3/C vdd NAND2X1
XNAND2X1_15 AND2X2_7/B AND2X2_7/A gnd NOR2X1_11/B vdd NAND2X1
XFILL_7_1 gnd vdd FILL
XNAND3X1_1 INVX2_8/Y INVX2_3/Y NAND3X1_1/C gnd AOI21X1_2/A vdd NAND3X1
XNAND2X1_27 A[2] INVX1_9/Y gnd NAND2X1_27/Y vdd NAND2X1
XFILL_1_1_0 gnd vdd FILL
XAOI22X1_6 INVX2_13/A AND2X2_2/Y A[2] INVX1_14/A gnd AOI22X1_6/Y vdd AOI22X1
XNAND2X1_16 NOR2X1_11/A NOR2X1_11/B gnd INVX1_7/A vdd NAND2X1
XFILL_6_0_0 gnd vdd FILL
XXOR2X1_1 B[1] A[1] gnd XOR2X1_1/Y vdd XOR2X1
XFILL_7_2 gnd vdd FILL
XNAND3X1_2 NAND3X1_2/A NAND2X1_1/Y NAND3X1_2/C gnd NAND3X1_2/Y vdd NAND3X1
XNAND2X1_17 INVX2_8/A AOI21X1_1/B gnd OAI21X1_6/C vdd NAND2X1
XNAND2X1_28 AND2X2_7/Y AOI21X1_8/B gnd INVX1_13/A vdd NAND2X1
XAOI22X1_7 AND2X2_7/A NOR2X1_1/B AND2X2_7/Y INVX2_12/A gnd AOI22X1_7/Y vdd AOI22X1
XFILL_1_1_1 gnd vdd FILL
XFILL_6_0_1 gnd vdd FILL
XXOR2X1_2 A[3] B[3] gnd XOR2X1_2/Y vdd XOR2X1
XFILL_7_3 gnd vdd FILL
XNAND2X1_18 A[6] B[6] gnd NAND3X1_7/B vdd NAND2X1
XNAND2X1_29 INVX4_2/Y AOI21X1_8/Y gnd NAND3X1_5/B vdd NAND2X1
XAOI22X1_8 AND2X2_1/A NOR2X1_1/B AND2X2_1/Y INVX2_12/A gnd AOI22X1_8/Y vdd AOI22X1
XNAND3X1_3 NAND3X1_3/A INVX1_15/A NAND3X1_3/C gnd NAND3X1_4/A vdd NAND3X1
XXOR2X1_3 A[2] B[2] gnd XOR2X1_3/Y vdd XOR2X1
XFILL_4_1_0 gnd vdd FILL
XINVX4_1 A[4] gnd INVX4_1/Y vdd INVX4
XOAI21X1_1 A[7] B[7] NOR2X1_1/B gnd NAND3X1_2/A vdd OAI21X1
XNAND2X1_19 A[0] B[0] gnd INVX2_9/A vdd NAND2X1
XAOI22X1_9 INVX1_14/A A[5] A[7] INVX4_3/A gnd AOI22X1_9/Y vdd AOI22X1
XNAND3X1_4 NAND3X1_4/A NAND3X1_4/B NAND3X1_4/C gnd BUFX2_3/A vdd NAND3X1
XINVX4_2 INVX4_2/A gnd INVX4_2/Y vdd INVX4
XFILL_4_1_1 gnd vdd FILL
XNAND3X1_5 INVX1_15/A NAND3X1_5/B NAND3X1_7/C gnd NAND3X1_5/Y vdd NAND3X1
XOAI21X1_2 INVX2_1/Y ALU_Sel[0] OR2X2_1/B gnd NOR2X1_1/A vdd OAI21X1
XINVX4_3 INVX4_3/A gnd INVX4_3/Y vdd INVX4
XNAND3X1_6 NAND3X1_5/Y NOR2X1_27/Y NAND3X1_6/C gnd BUFX2_7/A vdd NAND3X1
XOAI21X1_3 AND2X2_1/Y INVX1_3/Y INVX1_4/Y gnd INVX1_18/A vdd OAI21X1
XBUFX2_1 BUFX2_1/A gnd ALU_Out[0] vdd BUFX2
XNAND3X1_7 INVX2_8/A NAND3X1_7/B NAND3X1_7/C gnd NAND3X1_7/Y vdd NAND3X1
XINVX4_4 INVX4_4/A gnd INVX4_4/Y vdd INVX4
XINVX2_1 ALU_Sel[1] gnd INVX2_1/Y vdd INVX2
XAOI21X1_1 INVX2_8/A AOI21X1_1/B INVX4_4/Y gnd AOI21X1_1/Y vdd AOI21X1
XFILL_3_1 gnd vdd FILL
XOAI21X1_4 OAI21X1_4/A AOI21X1_3/Y OAI21X1_4/C gnd AOI21X1_5/B vdd OAI21X1
XAOI21X1_2 AOI21X1_2/A AOI21X1_1/Y NAND3X1_2/Y gnd NAND2X1_2/B vdd AOI21X1
XINVX2_2 A[6] gnd INVX2_2/Y vdd INVX2
XNAND3X1_8 INVX1_15/A NAND3X1_7/Y AOI22X1_2/A gnd NAND3X1_8/Y vdd NAND3X1
XBUFX2_2 BUFX2_2/A gnd ALU_Out[1] vdd BUFX2
XOAI21X1_5 AOI21X1_5/Y INVX4_2/A INVX2_3/Y gnd AOI21X1_1/B vdd OAI21X1
XAOI21X1_10 INVX2_11/Y NAND2X1_9/Y INVX4_4/Y gnd OAI21X1_19/C vdd AOI21X1
XFILL_3_2 gnd vdd FILL
XBUFX2_3 BUFX2_3/A gnd ALU_Out[2] vdd BUFX2
XOAI21X1_6 INVX1_1/Y B[7] OAI21X1_6/C gnd OAI21X1_6/Y vdd OAI21X1
XNOR2X1_1 NOR2X1_1/A NOR2X1_1/B gnd NOR2X1_1/Y vdd NOR2X1
XINVX2_3 INVX2_3/A gnd INVX2_3/Y vdd INVX2
XAOI21X1_3 AOI21X1_9/B NAND2X1_9/Y NOR2X1_6/Y gnd AOI21X1_3/Y vdd AOI21X1
XAOI21X1_11 AOI21X1_3/Y XOR2X1_3/Y INVX4_4/Y gnd OAI21X1_22/C vdd AOI21X1
XFILL_2_0_0 gnd vdd FILL
XNOR2X1_2 ALU_Sel[2] NOR2X1_2/B gnd INVX4_4/A vdd NOR2X1
XBUFX2_4 BUFX2_4/A gnd ALU_Out[3] vdd BUFX2
XAOI21X1_4 AOI21X1_4/A NOR2X1_8/Y NOR2X1_7/Y gnd OAI21X1_4/C vdd AOI21X1
XINVX2_4 A[5] gnd INVX2_4/Y vdd INVX2
XAOI21X1_12 INVX1_12/Y NAND3X1_3/A XOR2X1_2/Y gnd OAI21X1_28/B vdd AOI21X1
XOAI21X1_7 NOR2X1_11/A AND2X2_7/B AND2X2_1/B gnd OAI21X1_7/Y vdd OAI21X1
XFILL_1_1 gnd vdd FILL
XFILL_2_0_1 gnd vdd FILL
XNOR2X1_3 B[6] INVX2_2/Y gnd INVX2_3/A vdd NOR2X1
XINVX2_5 A[1] gnd INVX2_5/Y vdd INVX2
XOAI21X1_8 AOI21X1_6/Y OAI21X1_8/B AOI21X1_7/Y gnd AOI21X1_8/B vdd OAI21X1
XBUFX2_5 BUFX2_5/A gnd ALU_Out[4] vdd BUFX2
XAOI21X1_13 NOR2X1_11/B AOI21X1_5/B INVX4_4/Y gnd OAI21X1_34/C vdd AOI21X1
XAOI21X1_5 INVX1_7/Y AOI21X1_5/B INVX1_18/A gnd AOI21X1_5/Y vdd AOI21X1
XAOI21X1_6 INVX2_9/Y XOR2X1_1/Y NOR2X1_9/Y gnd AOI21X1_6/Y vdd AOI21X1
XNAND2X1_1 A[6] INVX1_14/A gnd NAND2X1_1/Y vdd NAND2X1
XINVX2_6 A[3] gnd INVX2_6/Y vdd INVX2
XFILL_0_1_0 gnd vdd FILL
XBUFX2_6 BUFX2_6/A gnd ALU_Out[5] vdd BUFX2
XOAI21X1_9 AOI21X1_8/Y INVX4_2/Y NAND3X1_7/B gnd OAI21X1_9/Y vdd OAI21X1
XNOR2X1_4 B[4] INVX4_1/Y gnd INVX1_3/A vdd NOR2X1
XAOI21X1_14 NOR2X1_25/Y AOI21X1_14/B AOI21X1_14/C gnd OAI21X1_45/A vdd AOI21X1
XFILL_5_0_0 gnd vdd FILL
XNOR2X1_5 B[5] INVX2_4/Y gnd INVX1_4/A vdd NOR2X1
XNAND2X1_2 NAND3X1_8/Y NAND2X1_2/B gnd BUFX2_8/A vdd NAND2X1
XBUFX2_7 BUFX2_7/A gnd ALU_Out[6] vdd BUFX2
XAOI21X1_7 INVX1_12/A XOR2X1_2/Y AND2X2_2/Y gnd AOI21X1_7/Y vdd AOI21X1
XFILL_0_1_1 gnd vdd FILL
XAOI21X1_15 INVX4_4/A XNOR2X1_6/Y OR2X2_2/Y gnd OAI21X1_42/C vdd AOI21X1
XINVX2_7 A[2] gnd INVX2_7/Y vdd INVX2
XFILL_5_0_1 gnd vdd FILL
XBUFX2_8 BUFX2_8/A gnd ALU_Out[7] vdd BUFX2
XINVX2_8 INVX2_8/A gnd INVX2_8/Y vdd INVX2
XNAND2X1_3 ALU_Sel[0] INVX2_1/Y gnd NOR2X1_2/B vdd NAND2X1
XAOI21X1_8 INVX1_17/A AOI21X1_8/B OAI21X1_7/Y gnd AOI21X1_8/Y vdd AOI21X1
XNOR2X1_6 B[1] INVX2_5/Y gnd NOR2X1_6/Y vdd NOR2X1
XAOI21X1_16 AOI21X1_7/Y OAI21X1_43/Y INVX1_17/Y gnd AOI21X1_16/Y vdd AOI21X1
XFILL_3_1_0 gnd vdd FILL
XBUFX2_9 BUFX2_9/A gnd CarryOut vdd BUFX2
XINVX2_9 INVX2_9/A gnd INVX2_9/Y vdd INVX2
XNAND2X1_4 B[6] INVX2_2/Y gnd NAND2X1_4/Y vdd NAND2X1
XAOI21X1_9 AOI21X1_9/A AOI21X1_9/B INVX2_9/A gnd AOI21X1_9/Y vdd AOI21X1
XAOI21X1_17 INVX4_2/Y NAND2X1_30/B INVX4_4/Y gnd OAI21X1_46/C vdd AOI21X1
XNOR2X1_7 B[3] INVX2_6/Y gnd NOR2X1_7/Y vdd NOR2X1
XNAND2X1_5 NAND2X1_4/Y INVX2_3/Y gnd INVX4_2/A vdd NAND2X1
XFILL_3_1_1 gnd vdd FILL
XNOR2X1_8 B[2] INVX2_7/Y gnd NOR2X1_8/Y vdd NOR2X1
XINVX1_10 B[0] gnd INVX1_10/Y vdd INVX1
XNOR2X1_9 INVX1_8/Y INVX2_5/Y gnd NOR2X1_9/Y vdd NOR2X1
XNAND2X1_6 A[5] B[5] gnd AND2X2_1/B vdd NAND2X1
XNAND2X1_7 INVX2_4/Y INVX1_2/Y gnd AND2X2_1/A vdd NAND2X1
XFILL_6_1_0 gnd vdd FILL
XINVX1_11 ALU_Sel[0] gnd INVX1_11/Y vdd INVX1
XFILL_6_1_1 gnd vdd FILL
XNAND2X1_8 B[1] INVX2_5/Y gnd AOI21X1_9/B vdd NAND2X1
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XNOR2X1_20 NOR2X1_20/A NOR2X1_20/B gnd NAND3X1_4/C vdd NOR2X1
XOAI21X1_40 OAI21X1_45/A AND2X2_7/Y INVX1_3/Y gnd XNOR2X1_6/A vdd OAI21X1
XNOR2X1_10 INVX2_7/Y INVX1_9/Y gnd INVX1_12/A vdd NOR2X1
XNOR2X1_21 NOR2X1_26/A NOR2X1_21/B gnd NOR2X1_21/Y vdd NOR2X1
XNAND2X1_9 B[0] INVX1_5/Y gnd NAND2X1_9/Y vdd NAND2X1
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XFILL_6_1 gnd vdd FILL
XOAI21X1_30 INVX2_12/Y NOR2X1_26/A OAI21X1_30/C gnd NOR2X1_22/A vdd OAI21X1
XOAI21X1_41 AND2X2_1/B INVX2_13/Y AOI22X1_8/Y gnd OR2X2_2/A vdd OAI21X1
XFILL_1_0_0 gnd vdd FILL
XNOR2X1_22 NOR2X1_22/A NOR2X1_22/B gnd AND2X2_6/B vdd NOR2X1
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XNOR2X1_11 NOR2X1_11/A NOR2X1_11/B gnd INVX1_17/A vdd NOR2X1
XOAI21X1_20 AOI21X1_9/Y OAI21X1_20/B AND2X2_5/Y gnd BUFX2_2/A vdd OAI21X1
XOAI21X1_31 INVX4_1/Y INVX4_3/Y AOI22X1_6/Y gnd NOR2X1_22/B vdd OAI21X1
XOAI21X1_42 XNOR2X1_5/Y INVX1_15/Y OAI21X1_42/C gnd BUFX2_6/A vdd OAI21X1
XFILL_1_0_1 gnd vdd FILL
XNOR2X1_12 AND2X2_3/Y INVX4_4/A gnd AOI22X1_2/B vdd NOR2X1
XNOR2X1_23 NOR2X1_23/A NOR2X1_23/B gnd AND2X2_8/B vdd NOR2X1
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XOAI21X1_10 NOR2X1_2/B ALU_Sel[2] NOR2X1_16/B gnd OAI21X1_10/Y vdd OAI21X1
XOAI21X1_43 AOI21X1_9/Y NOR2X1_9/Y NOR2X1_26/Y gnd OAI21X1_43/Y vdd OAI21X1
XOAI21X1_21 AOI21X1_9/Y NOR2X1_9/Y XOR2X1_3/Y gnd NAND3X1_3/A vdd OAI21X1
XOAI21X1_32 INVX4_4/Y XNOR2X1_4/Y AND2X2_6/Y gnd BUFX2_4/A vdd OAI21X1
XNOR2X1_24 A[0] INVX1_10/Y gnd NOR2X1_24/Y vdd NOR2X1
XNOR2X1_13 ALU_Sel[2] NOR2X1_14/B gnd INVX2_13/A vdd NOR2X1
XINVX1_16 NOR2X1_7/Y gnd INVX1_16/Y vdd INVX1
XOAI21X1_11 INVX1_5/Y INVX1_10/Y OAI21X1_10/Y gnd OAI21X1_11/Y vdd OAI21X1
XOAI21X1_44 AOI21X1_16/Y OAI21X1_7/Y INVX4_2/A gnd NAND3X1_7/C vdd OAI21X1
XOAI21X1_22 AOI21X1_3/Y XOR2X1_3/Y OAI21X1_22/C gnd NAND3X1_4/B vdd OAI21X1
XOAI21X1_33 AOI21X1_8/B AND2X2_7/Y INVX1_15/A gnd OAI21X1_36/B vdd OAI21X1
XFILL_4_0_0 gnd vdd FILL
XFILL_4_1 gnd vdd FILL
XNOR2X1_14 OR2X2_1/B NOR2X1_14/B gnd INVX4_3/A vdd NOR2X1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XNOR2X1_25 XOR2X1_2/Y XOR2X1_3/Y gnd NOR2X1_25/Y vdd NOR2X1
XOAI21X1_12 ALU_Sel[2] OR2X2_1/A OAI21X1_11/Y gnd OAI21X1_13/C vdd OAI21X1
XFILL_4_0_1 gnd vdd FILL
XOAI21X1_45 OAI21X1_45/A INVX1_7/A INVX1_18/Y gnd NAND2X1_30/B vdd OAI21X1
XOAI21X1_23 A[2] B[2] NOR2X1_1/B gnd OAI21X1_24/C vdd OAI21X1
XOAI21X1_34 AOI21X1_5/B NOR2X1_11/B OAI21X1_34/C gnd AND2X2_8/A vdd OAI21X1
XNOR2X1_15 ALU_Sel[2] NOR2X1_16/B gnd INVX1_15/A vdd NOR2X1
XNOR2X1_26 NOR2X1_26/A NOR2X1_26/B gnd NOR2X1_26/Y vdd NOR2X1
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XOAI21X1_13 A[0] B[0] OAI21X1_13/C gnd AND2X2_4/A vdd OAI21X1
XOAI21X1_46 INVX4_2/Y NAND2X1_30/B OAI21X1_46/C gnd NAND3X1_6/C vdd OAI21X1
XOAI21X1_35 AND2X2_7/B INVX2_13/Y AOI22X1_7/Y gnd NOR2X1_23/B vdd OAI21X1
XOAI21X1_24 INVX2_12/Y NOR2X1_26/B OAI21X1_24/C gnd NOR2X1_20/A vdd OAI21X1
XNOR2X1_16 OR2X2_1/B NOR2X1_16/B gnd INVX2_12/A vdd NOR2X1
XNOR2X1_27 NOR2X1_27/A NOR2X1_27/B gnd NOR2X1_27/Y vdd NOR2X1
XFILL_2_1_0 gnd vdd FILL
XOAI21X1_14 OAI21X1_6/Y OR2X2_1/Y AND2X2_4/Y gnd BUFX2_1/A vdd OAI21X1
XOAI21X1_47 A[6] B[6] NOR2X1_1/B gnd OAI21X1_48/C vdd OAI21X1
XOAI21X1_25 INVX2_6/Y INVX4_3/Y AOI22X1_5/Y gnd NOR2X1_20/B vdd OAI21X1
XOAI21X1_36 INVX1_13/Y OAI21X1_36/B AND2X2_8/Y gnd BUFX2_5/A vdd OAI21X1
XXNOR2X1_1 A[7] B[7] gnd INVX2_8/A vdd XNOR2X1
XINVX1_1 A[7] gnd INVX1_1/Y vdd INVX1
XNOR2X1_17 ALU_Sel[2] OR2X2_1/A gnd NOR2X1_1/B vdd NOR2X1
XAND2X2_1 AND2X2_1/A AND2X2_1/B gnd AND2X2_1/Y vdd AND2X2
XFILL_2_1 gnd vdd FILL
XFILL_2_1_1 gnd vdd FILL
XOAI21X1_15 XOR2X1_1/Y INVX2_9/Y INVX1_15/A gnd OAI21X1_20/B vdd OAI21X1
XOAI21X1_48 INVX4_2/Y INVX2_12/Y OAI21X1_48/C gnd NOR2X1_27/B vdd OAI21X1
XOAI21X1_26 AOI21X1_3/Y XOR2X1_3/Y NAND2X1_27/Y gnd XNOR2X1_4/A vdd OAI21X1
XOAI21X1_37 INVX4_1/Y INVX1_6/Y INVX1_13/A gnd XNOR2X1_5/A vdd OAI21X1
XINVX1_2 B[5] gnd INVX1_2/Y vdd INVX1
XXNOR2X1_2 A[3] B[3] gnd NOR2X1_26/A vdd XNOR2X1
XAND2X2_2 A[3] B[3] gnd AND2X2_2/Y vdd AND2X2
XNOR2X1_18 OR2X2_1/B NOR2X1_2/B gnd INVX1_14/A vdd NOR2X1
XOAI21X1_16 B[1] A[1] NOR2X1_1/B gnd OAI21X1_17/C vdd OAI21X1
XOAI21X1_38 XOR2X1_1/Y NOR2X1_24/Y AOI21X1_9/A gnd AOI21X1_14/B vdd OAI21X1
XOAI21X1_49 NAND3X1_7/B INVX2_13/Y AOI22X1_9/Y gnd NOR2X1_27/A vdd OAI21X1
XOAI21X1_27 AOI21X1_6/Y NOR2X1_26/B INVX1_12/Y gnd NOR2X1_21/B vdd OAI21X1
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XXNOR2X1_3 A[2] B[2] gnd NOR2X1_26/B vdd XNOR2X1
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XAND2X2_3 A[7] B[7] gnd AND2X2_3/Y vdd AND2X2
XFILL_5_1_0 gnd vdd FILL
XNOR2X1_19 NOR2X1_19/A NOR2X1_19/B gnd AND2X2_5/A vdd NOR2X1
XNAND2X1_30 INVX4_2/Y NAND2X1_30/B gnd NAND3X1_1/C vdd NAND2X1
XOAI22X1_1 INVX1_14/Y INVX2_6/Y INVX2_4/Y INVX4_3/Y gnd NOR2X1_23/A vdd OAI22X1
XINVX2_10 ALU_Sel[2] gnd OR2X2_1/B vdd INVX2
XOAI21X1_17 INVX2_12/Y INVX2_11/Y OAI21X1_17/C gnd NOR2X1_19/A vdd OAI21X1
XOAI21X1_28 NOR2X1_21/Y OAI21X1_28/B INVX1_15/A gnd AND2X2_6/A vdd OAI21X1
XOAI21X1_39 XOR2X1_2/Y NAND2X1_27/Y INVX1_16/Y gnd AOI21X1_14/C vdd OAI21X1
XFILL_5_1_1 gnd vdd FILL
XXNOR2X1_4 XNOR2X1_4/A NOR2X1_26/A gnd XNOR2X1_4/Y vdd XNOR2X1
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XAND2X2_4 AND2X2_4/A AND2X2_4/B gnd AND2X2_4/Y vdd AND2X2
XNAND2X1_20 XOR2X1_2/Y XOR2X1_3/Y gnd OAI21X1_8/B vdd NAND2X1
XOAI21X1_18 INVX2_7/Y INVX4_3/Y AOI22X1_4/Y gnd NOR2X1_19/B vdd OAI21X1
XINVX2_11 XOR2X1_1/Y gnd INVX2_11/Y vdd INVX2
XOAI21X1_29 A[3] B[3] NOR2X1_1/B gnd OAI21X1_30/C vdd OAI21X1
XOAI22X1_2 INVX2_2/Y INVX4_3/Y INVX1_14/Y INVX4_1/Y gnd OR2X2_2/B vdd OAI22X1
XINVX1_5 A[0] gnd INVX1_5/Y vdd INVX1
XXNOR2X1_5 XNOR2X1_5/A AND2X2_1/Y gnd XNOR2X1_5/Y vdd XNOR2X1
.ends

