* NGSPICE file created from ALU.ext - technology: scmos

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

.subckt ALU vdd gnd A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] B[0] B[1] B[2] B[3] B[4]
+ B[5] B[6] B[7] opcode[0] opcode[1] opcode[2] opcode[3] result[0] result[1] result[2]
+ result[3] result[4] result[5] result[6] result[7] overflow negative zero
XAND2X2_5 B[3] A[3] gnd AND2X2_5/Y vdd AND2X2
XNAND2X1_21 A[0] B[0] gnd OAI21X1_2/B vdd NAND2X1
XOAI22X1_3 A[0] INVX1_16/Y AND2X2_3/Y NOR2X1_41/A gnd OAI22X1_3/Y vdd OAI22X1
XNAND2X1_32 AOI22X1_2/D OR2X2_4/Y gnd NOR2X1_43/B vdd NAND2X1
XNAND2X1_10 B[4] A[4] gnd INVX1_4/A vdd NAND2X1
XINVX2_12 A[2] gnd OR2X2_2/A vdd INVX2
XOAI21X1_19 INVX2_6/A AND2X2_2/B INVX2_1/A gnd NOR2X1_9/A vdd OAI21X1
XOR2X2_4 A[1] B[1] gnd OR2X2_4/Y vdd OR2X2
XFILL_0_0_0 gnd vdd FILL
XINVX1_6 INVX1_6/A gnd BUFX2_8/A vdd INVX1
XNAND2X1_22 opcode[0] NOR2X1_2/B gnd NOR2X1_38/A vdd NAND2X1
XAND2X2_6 A[0] B[0] gnd AND2X2_6/Y vdd AND2X2
XNAND2X1_33 OAI22X1_3/Y INVX2_1/A gnd OAI21X1_51/A vdd NAND2X1
XAOI22X1_1 OR2X2_2/A NOR2X1_38/Y INVX2_5/A XOR2X1_1/Y gnd OAI21X1_4/C vdd AOI22X1
XNAND2X1_11 INVX2_8/Y INVX2_4/Y gnd AOI22X1_6/B vdd NAND2X1
XINVX2_13 A[1] gnd OR2X2_3/A vdd INVX2
XOAI22X1_4 NOR2X1_5/A NOR2X1_26/Y AND2X2_5/Y OAI22X1_4/D gnd OAI22X1_4/Y vdd OAI22X1
XOR2X2_5 B[2] A[2] gnd OR2X2_5/Y vdd OR2X2
XFILL_0_0_1 gnd vdd FILL
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XNAND2X1_23 opcode[1] INVX1_18/Y gnd NOR2X1_36/A vdd NAND2X1
XAOI22X1_10 INVX2_10/Y NOR2X1_38/Y INVX2_19/A NOR2X1_20/B gnd AOI22X1_10/Y vdd AOI22X1
XAOI22X1_2 INVX2_15/Y B[0] OR2X2_4/Y AOI22X1_2/D gnd AOI22X1_2/Y vdd AOI22X1
XNAND2X1_12 INVX2_6/Y INVX2_2/Y gnd AOI21X1_7/C vdd NAND2X1
XNAND2X1_34 B[2] A[2] gnd OAI21X1_8/A vdd NAND2X1
XINVX2_14 INVX2_14/A gnd INVX2_14/Y vdd INVX2
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XAOI22X1_3 INVX1_14/Y NOR2X1_38/Y INVX2_5/A XOR2X1_3/Y gnd NAND3X1_4/B vdd AOI22X1
XNAND2X1_24 opcode[2] INVX1_19/Y gnd NOR2X1_42/A vdd NAND2X1
XAOI22X1_11 INVX2_15/Y INVX1_16/Y AOI22X1_11/C INVX2_17/Y gnd NOR2X1_39/B vdd AOI22X1
XINVX2_15 A[0] gnd INVX2_15/Y vdd INVX2
XNAND2X1_13 INVX2_6/A INVX2_2/A gnd INVX1_8/A vdd NAND2X1
XNOR3X1_1 NOR3X1_1/A NOR3X1_1/B NOR3X1_1/C gnd NOR3X1_1/Y vdd NOR3X1
XFILL_3_0_0 gnd vdd FILL
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XNAND2X1_25 A[0] NOR2X1_40/Y gnd NAND2X1_25/Y vdd NAND2X1
XAOI22X1_12 INVX1_3/A A[1] INVX2_15/Y NOR2X1_38/Y gnd AOI22X1_12/Y vdd AOI22X1
XNAND2X1_14 B[5] A[5] gnd NAND2X1_14/Y vdd NAND2X1
XNOR3X1_2 NOR3X1_2/A NOR3X1_2/B NOR3X1_2/C gnd NOR3X1_2/Y vdd NOR3X1
XAOI22X1_4 INVX2_17/A OR2X2_1/Y AND2X2_5/Y INVX2_19/A gnd AOI22X1_4/Y vdd AOI22X1
XINVX2_16 INVX2_16/A gnd INVX2_16/Y vdd INVX2
XFILL_3_0_1 gnd vdd FILL
XINVX2_17 INVX2_17/A gnd INVX2_17/Y vdd INVX2
XNAND2X1_15 INVX2_11/Y NOR2X1_38/Y gnd OAI21X1_33/C vdd NAND2X1
XNAND2X1_26 OR2X2_3/A NOR2X1_38/Y gnd NAND2X1_26/Y vdd NAND2X1
XAOI22X1_5 INVX1_3/A A[4] A[2] NOR2X1_40/Y gnd NAND3X1_4/A vdd AOI22X1
XNOR3X1_3 NOR3X1_3/A NOR3X1_3/B NOR3X1_3/C gnd NOR3X1_3/Y vdd NOR3X1
XFILL_7_1 gnd vdd FILL
XNAND2X1_16 NOR2X1_15/Y NAND3X1_8/Y gnd AOI21X1_16/C vdd NAND2X1
XNAND2X1_27 NOR2X1_41/Y INVX2_5/A gnd NAND2X1_27/Y vdd NAND2X1
XNAND3X1_1 NAND3X1_1/A NAND3X1_1/B OAI21X1_5/Y gnd NOR3X1_1/A vdd NAND3X1
XNOR3X1_4 BUFX2_3/A BUFX2_6/A NOR3X1_4/C gnd NOR3X1_4/Y vdd NOR3X1
XAOI22X1_6 INVX2_17/A AOI22X1_6/B INVX1_4/Y INVX2_19/A gnd AOI22X1_6/Y vdd AOI22X1
XFILL_1_1_0 gnd vdd FILL
XINVX2_18 INVX2_18/A gnd INVX2_18/Y vdd INVX2
XFILL_6_0_0 gnd vdd FILL
XXOR2X1_1 B[2] A[2] gnd XOR2X1_1/Y vdd XOR2X1
XFILL_7_2 gnd vdd FILL
XNAND3X1_2 OR2X2_2/Y XOR2X1_3/Y OAI21X1_6/Y gnd NAND3X1_2/Y vdd NAND3X1
XNAND2X1_17 NAND3X1_7/Y NAND2X1_17/B gnd BUFX2_1/A vdd NAND2X1
XNAND2X1_28 AND2X2_3/Y INVX2_19/A gnd NAND3X1_16/C vdd NAND2X1
XNOR3X1_5 BUFX2_9/A BUFX2_1/A NOR3X1_5/C gnd NOR3X1_5/Y vdd NOR3X1
XFILL_1_1_1 gnd vdd FILL
XAOI22X1_7 NOR2X1_38/Y INVX2_4/Y A[3] NOR2X1_40/Y gnd AOI22X1_7/Y vdd AOI22X1
XFILL_6_0_1 gnd vdd FILL
XINVX2_19 INVX2_19/A gnd INVX2_19/Y vdd INVX2
XXOR2X1_2 B[5] A[5] gnd INVX2_6/A vdd XOR2X1
XNOR3X1_6 NOR3X1_6/A A[7] NOR3X1_6/C gnd NOR3X1_6/Y vdd NOR3X1
XNAND2X1_29 A[2] INVX1_3/A gnd NAND3X1_16/A vdd NAND2X1
XNAND2X1_18 A[5] INVX1_11/Y gnd OAI21X1_42/C vdd NAND2X1
XAOI22X1_8 OR2X2_5/Y OAI21X1_8/A NAND2X1_6/Y OR2X2_1/Y gnd AOI22X1_8/Y vdd AOI22X1
XNAND3X1_3 XOR2X1_1/Y XOR2X1_3/Y AOI21X1_2/B gnd AOI21X1_4/A vdd NAND3X1
XXOR2X1_3 B[3] A[3] gnd XOR2X1_3/Y vdd XOR2X1
XINVX4_1 INVX4_1/A gnd INVX4_1/Y vdd INVX4
XFILL_4_1_0 gnd vdd FILL
XNOR3X1_7 NOR3X1_6/Y NOR3X1_7/B NOR3X1_7/C gnd BUFX2_2/A vdd NOR3X1
XAOI22X1_9 INVX1_3/A A[6] INVX1_2/Y NOR2X1_38/Y gnd AOI22X1_9/Y vdd AOI22X1
XNAND3X1_4 NAND3X1_4/A NAND3X1_4/B AOI22X1_4/Y gnd AOI21X1_4/C vdd NAND3X1
XNAND2X1_19 A[4] INVX2_8/Y gnd AND2X2_2/B vdd NAND2X1
XOAI21X1_1 OAI21X1_1/A NOR3X1_3/A NOR2X1_1/Y gnd NAND3X1_9/A vdd OAI21X1
XXOR2X1_4 B[4] A[4] gnd INVX2_2/A vdd XOR2X1
XNAND3X1_5 NAND3X1_5/A NAND3X1_5/B NAND3X1_5/C gnd BUFX2_9/A vdd NAND3X1
XFILL_4_1_1 gnd vdd FILL
XNOR3X1_8 NOR3X1_8/A NOR3X1_8/B NOR3X1_8/C gnd INVX1_20/A vdd NOR3X1
XOAI21X1_2 NOR2X1_41/A OAI21X1_2/B AOI22X1_2/D gnd AOI21X1_2/B vdd OAI21X1
XNAND3X1_6 INVX4_1/A INVX1_10/Y NAND3X1_6/C gnd NAND3X1_7/B vdd NAND3X1
XOAI21X1_3 XOR2X1_1/Y AOI21X1_2/B INVX2_7/A gnd AOI21X1_2/C vdd OAI21X1
XFILL_7_1_0 gnd vdd FILL
XBUFX2_1 BUFX2_1/A gnd negative vdd BUFX2
XNAND3X1_7 INVX2_1/A NAND3X1_7/B NAND3X1_7/C gnd NAND3X1_7/Y vdd NAND3X1
XAOI21X1_20 A[7] INVX1_12/Y opcode[2] gnd NAND3X1_13/C vdd AOI21X1
XINVX2_1 INVX2_1/A gnd INVX2_1/Y vdd INVX2
XAOI21X1_1 OR2X2_3/Y OAI22X1_3/Y XOR2X1_1/Y gnd NOR2X1_1/B vdd AOI21X1
XOAI21X1_4 OR2X2_3/A NAND2X1_2/Y OAI21X1_4/C gnd NOR3X1_1/C vdd OAI21X1
XFILL_3_1 gnd vdd FILL
XFILL_7_1_1 gnd vdd FILL
XBUFX2_2 BUFX2_2/A gnd overflow vdd BUFX2
XNAND3X1_8 INVX1_9/Y NAND3X1_8/B NAND3X1_8/C gnd NAND3X1_8/Y vdd NAND3X1
XAOI21X1_2 XOR2X1_1/Y AOI21X1_2/B AOI21X1_2/C gnd NOR3X1_1/B vdd AOI21X1
XINVX2_2 INVX2_2/A gnd INVX2_2/Y vdd INVX2
XAOI21X1_21 INVX1_10/A INVX4_1/Y AOI21X1_21/C gnd OAI21X1_44/C vdd AOI21X1
XOAI21X1_5 B[2] A[2] INVX2_17/A gnd OAI21X1_5/Y vdd OAI21X1
XAOI21X1_10 AOI21X1_10/A NOR2X1_9/Y OAI21X1_25/Y gnd INVX1_6/A vdd AOI21X1
XBUFX2_3 BUFX2_3/A gnd result[0] vdd BUFX2
XNAND3X1_9 NAND3X1_9/A INVX1_20/A NOR3X1_1/Y gnd NOR3X1_4/C vdd NAND3X1
XBUFX2_10 BUFX2_1/A gnd result[7] vdd BUFX2
XAOI21X1_11 INVX2_9/Y OAI21X1_27/Y INVX2_14/A gnd NOR2X1_11/B vdd AOI21X1
XAOI21X1_22 OR2X2_3/Y OAI22X1_3/Y OAI22X1_4/Y gnd NOR2X1_28/B vdd AOI21X1
XAOI21X1_3 NAND2X1_9/Y NOR2X1_5/Y OAI21X1_8/Y gnd AOI21X1_3/Y vdd AOI21X1
XINVX2_3 INVX2_3/A gnd INVX2_3/Y vdd INVX2
XOAI21X1_6 AOI22X1_2/Y NOR2X1_3/Y NOR3X1_3/A gnd OAI21X1_6/Y vdd OAI21X1
XNOR2X1_1 INVX2_1/Y NOR2X1_1/B gnd NOR2X1_1/Y vdd NOR2X1
XFILL_2_0_0 gnd vdd FILL
XNOR2X1_2 opcode[0] NOR2X1_2/B gnd NOR2X1_2/Y vdd NOR2X1
XBUFX2_4 BUFX2_4/A gnd result[1] vdd BUFX2
XBUFX2_11 NOR3X1_5/Y gnd zero vdd BUFX2
XAOI21X1_4 AOI21X1_4/A AOI21X1_3/Y AOI21X1_4/C gnd AOI21X1_4/Y vdd AOI21X1
XINVX2_4 A[4] gnd INVX2_4/Y vdd INVX2
XAOI21X1_12 AND2X2_6/Y OR2X2_4/Y AND2X2_3/Y gnd NOR3X1_3/C vdd AOI21X1
XOAI21X1_7 NOR2X1_1/B NOR2X1_4/Y NOR3X1_3/B gnd OAI21X1_7/Y vdd OAI21X1
XFILL_1_1 gnd vdd FILL
XFILL_2_0_1 gnd vdd FILL
XINVX2_5 INVX2_5/A gnd INVX2_5/Y vdd INVX2
XAOI21X1_13 INVX1_7/Y OAI21X1_31/Y INVX2_14/Y gnd NOR2X1_12/B vdd AOI21X1
XNOR2X1_3 B[1] OR2X2_3/A gnd NOR2X1_3/Y vdd NOR2X1
XOAI21X1_8 OAI21X1_8/A NOR3X1_3/B INVX2_7/A gnd OAI21X1_8/Y vdd OAI21X1
XAOI21X1_5 NOR2X1_31/A INVX2_2/A AOI21X1_5/C gnd NOR2X1_8/A vdd AOI21X1
XBUFX2_5 BUFX2_5/A gnd result[2] vdd BUFX2
XFILL_1_2 gnd vdd FILL
XAOI21X1_6 NOR2X1_4/Y NOR3X1_3/B INVX1_15/A gnd AOI21X1_7/A vdd AOI21X1
XINVX2_6 INVX2_6/A gnd INVX2_6/Y vdd INVX2
XNAND2X1_1 OAI21X1_8/A OR2X2_5/Y gnd NOR3X1_3/A vdd NAND2X1
XBUFX2_6 BUFX2_6/A gnd result[3] vdd BUFX2
XFILL_0_1_0 gnd vdd FILL
XAOI21X1_14 A[5] NOR2X1_40/Y OAI21X1_33/Y gnd AOI21X1_14/Y vdd AOI21X1
XNOR2X1_4 B[2] OR2X2_2/A gnd NOR2X1_4/Y vdd NOR2X1
XOAI21X1_9 INVX2_1/Y OAI21X1_9/B AOI21X1_4/Y gnd BUFX2_6/A vdd OAI21X1
XFILL_5_0_0 gnd vdd FILL
XBUFX2_7 INVX1_5/Y gnd result[4] vdd BUFX2
XNAND2X1_2 NOR2X1_2/Y AND2X2_1/Y gnd NAND2X1_2/Y vdd NAND2X1
XINVX2_7 INVX2_7/A gnd INVX2_7/Y vdd INVX2
XNOR2X1_5 NOR2X1_5/A XOR2X1_3/Y gnd NOR2X1_5/Y vdd NOR2X1
XFILL_0_1_1 gnd vdd FILL
XAOI21X1_15 INVX1_1/Y AOI21X1_4/A INVX1_8/A gnd AOI21X1_15/Y vdd AOI21X1
XAOI21X1_7 AOI21X1_7/A AOI21X1_7/B AOI21X1_7/C gnd NOR2X1_9/B vdd AOI21X1
XFILL_5_0_1 gnd vdd FILL
XNAND2X1_3 NOR2X1_5/A INVX2_19/A gnd NAND3X1_1/B vdd NAND2X1
XINVX2_8 B[4] gnd INVX2_8/Y vdd INVX2
XAOI21X1_8 INVX2_2/A INVX2_3/A AOI21X1_8/C gnd AOI21X1_8/Y vdd AOI21X1
XBUFX2_8 BUFX2_8/A gnd result[5] vdd BUFX2
XAOI21X1_16 OAI21X1_38/Y NOR2X1_14/Y AOI21X1_16/C gnd NAND2X1_17/B vdd AOI21X1
XNOR2X1_6 INVX2_2/Y INVX2_3/Y gnd NOR2X1_6/Y vdd NOR2X1
XFILL_3_1_0 gnd vdd FILL
XAOI21X1_17 AOI21X1_17/A AOI21X1_17/B INVX2_1/Y gnd NOR3X1_6/A vdd AOI21X1
XBUFX2_9 BUFX2_9/A gnd result[6] vdd BUFX2
XINVX2_9 INVX2_9/A gnd INVX2_9/Y vdd INVX2
XAOI21X1_9 INVX1_4/Y INVX2_6/A INVX2_7/Y gnd AOI21X1_9/Y vdd AOI21X1
XNAND2X1_4 A[3] INVX1_3/A gnd NAND3X1_1/A vdd NAND2X1
XNOR2X1_7 NOR2X1_7/A NOR2X1_7/B gnd NOR2X1_7/Y vdd NOR2X1
XFILL_3_1_1 gnd vdd FILL
XNAND2X1_5 NAND3X1_9/A NOR3X1_1/Y gnd BUFX2_5/A vdd NAND2X1
XAOI21X1_18 INVX4_1/A INVX2_1/A NOR2X1_14/Y gnd NOR3X1_7/B vdd AOI21X1
XINVX1_20 INVX1_20/A gnd BUFX2_4/A vdd INVX1
XNOR2X1_8 NOR2X1_8/A NOR2X1_8/B gnd INVX1_5/A vdd NOR2X1
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XNOR2X1_40 NOR2X1_36/A NOR2X1_42/A gnd NOR2X1_40/Y vdd NOR2X1
XNOR2X1_9 NOR2X1_9/A NOR2X1_9/B gnd NOR2X1_9/Y vdd NOR2X1
XNAND2X1_6 B[3] A[3] gnd NAND2X1_6/Y vdd NAND2X1
XFILL_8_1 gnd vdd FILL
XAOI21X1_19 NAND3X1_7/Y NAND2X1_17/B INVX2_10/Y gnd NOR3X1_7/C vdd AOI21X1
XFILL_6_1_0 gnd vdd FILL
XNOR2X1_41 NOR2X1_41/A AND2X2_3/Y gnd NOR2X1_41/Y vdd NOR2X1
XNOR2X1_30 INVX2_6/A INVX2_2/A gnd NOR2X1_30/Y vdd NOR2X1
XNAND2X1_7 NAND2X1_6/Y OR2X2_1/Y gnd NOR3X1_3/B vdd NAND2X1
XINVX1_11 B[5] gnd INVX1_11/Y vdd INVX1
XOAI21X1_50 AND2X2_3/Y NOR2X1_41/A OAI21X1_2/B gnd OAI21X1_50/Y vdd OAI21X1
XFILL_6_1_1 gnd vdd FILL
XNOR2X1_20 NOR2X1_20/A NOR2X1_20/B gnd INVX4_1/A vdd NOR2X1
XINVX1_12 B[7] gnd INVX1_12/Y vdd INVX1
XNOR2X1_42 NOR2X1_42/A INVX2_18/Y gnd INVX2_5/A vdd NOR2X1
XNOR2X1_31 NOR2X1_31/A NOR2X1_31/B gnd NOR2X1_31/Y vdd NOR2X1
XNAND2X1_8 NAND3X1_2/Y OAI21X1_7/Y gnd OAI21X1_9/B vdd NAND2X1
XOAI21X1_40 NOR2X1_11/B INVX1_10/A INVX4_1/A gnd AOI21X1_17/B vdd OAI21X1
XOAI21X1_51 OAI21X1_51/A NOR2X1_43/Y NAND3X1_18/Y gnd NOR3X1_8/C vdd OAI21X1
XNOR2X1_32 opcode[3] opcode[2] gnd INVX2_16/A vdd NOR2X1
XNOR2X1_21 B[6] INVX2_11/Y gnd INVX1_10/A vdd NOR2X1
XNOR2X1_43 NOR2X1_43/A NOR2X1_43/B gnd NOR2X1_43/Y vdd NOR2X1
XNOR2X1_10 INVX2_4/Y NAND2X1_2/Y gnd NOR3X1_2/B vdd NOR2X1
XNAND3X1_10 INVX1_5/A INVX1_6/A NOR3X1_4/Y gnd NOR3X1_5/C vdd NAND3X1
XINVX1_13 B[6] gnd INVX1_13/Y vdd INVX1
XNAND2X1_9 XOR2X1_1/Y AOI21X1_2/B gnd NAND2X1_9/Y vdd NAND2X1
XOAI21X1_41 NOR2X1_12/B INVX1_9/A NOR2X1_14/Y gnd OAI21X1_41/Y vdd OAI21X1
XOAI21X1_30 INVX2_3/Y INVX1_8/A INVX1_7/Y gnd OAI21X1_30/Y vdd OAI21X1
XOAI21X1_52 OR2X2_3/A B[1] OAI22X1_3/Y gnd OAI21X1_1/A vdd OAI21X1
XFILL_1_0_0 gnd vdd FILL
XNAND3X1_11 INVX4_1/Y INVX1_10/Y NAND3X1_6/C gnd AOI21X1_17/A vdd NAND3X1
XNOR2X1_44 INVX2_18/Y INVX2_16/Y gnd INVX2_7/A vdd NOR2X1
XNOR2X1_33 NOR2X1_33/A INVX2_16/Y gnd INVX2_17/A vdd NOR2X1
XNOR2X1_22 INVX1_13/Y INVX2_11/Y gnd INVX1_9/A vdd NOR2X1
XNOR2X1_11 INVX2_1/Y NOR2X1_11/B gnd NOR2X1_11/Y vdd NOR2X1
XINVX1_14 A[3] gnd INVX1_14/Y vdd INVX1
XOAI21X1_42 INVX2_6/A AND2X2_2/B OAI21X1_42/C gnd INVX2_9/A vdd OAI21X1
XOAI21X1_31 NOR3X1_3/Y INVX1_1/A INVX1_8/Y gnd OAI21X1_31/Y vdd OAI21X1
XOAI21X1_20 INVX2_8/Y INVX2_4/Y INVX2_6/Y gnd AOI21X1_8/C vdd OAI21X1
XFILL_1_0_1 gnd vdd FILL
XNAND3X1_12 NOR2X1_15/Y NAND3X1_8/Y OAI21X1_41/Y gnd NOR3X1_6/C vdd NAND3X1
XNOR2X1_12 INVX2_7/Y NOR2X1_12/B gnd NOR2X1_12/Y vdd NOR2X1
XNOR2X1_34 NOR2X1_38/A INVX2_16/Y gnd INVX2_1/A vdd NOR2X1
XNOR2X1_23 B[6] A[6] gnd NOR2X1_23/Y vdd NOR2X1
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XOAI21X1_43 INVX1_9/A NOR2X1_23/Y INVX4_1/Y gnd OAI21X1_44/A vdd OAI21X1
XOAI21X1_32 INVX2_14/A OAI21X1_30/Y NOR2X1_12/Y gnd NAND3X1_5/C vdd OAI21X1
XOAI21X1_21 INVX2_3/Y INVX1_8/A AOI21X1_9/Y gnd OAI21X1_25/A vdd OAI21X1
XOAI21X1_10 NOR2X1_31/A INVX2_2/A INVX2_1/A gnd AOI21X1_5/C vdd OAI21X1
XNAND3X1_13 opcode[3] INVX2_18/A NAND3X1_13/C gnd AOI21X1_21/C vdd NAND3X1
XNOR2X1_35 opcode[3] INVX2_18/Y gnd NOR2X1_35/Y vdd NOR2X1
XNOR2X1_13 NOR2X1_13/A NOR2X1_13/B gnd NAND3X1_5/B vdd NOR2X1
XINVX1_16 B[0] gnd INVX1_16/Y vdd INVX1
XNOR2X1_24 B[3] INVX1_14/Y gnd INVX1_15/A vdd NOR2X1
XOAI21X1_44 OAI21X1_44/A INVX2_9/Y OAI21X1_44/C gnd OAI21X1_48/B vdd OAI21X1
XOAI21X1_33 INVX2_14/Y INVX2_5/Y OAI21X1_33/C gnd OAI21X1_33/Y vdd OAI21X1
XOAI21X1_22 INVX2_6/Y INVX2_5/Y AOI22X1_9/Y gnd NOR3X1_2/C vdd OAI21X1
XOAI21X1_11 OAI22X1_4/D OAI21X1_8/A NAND2X1_6/Y gnd INVX1_1/A vdd OAI21X1
XFILL_4_0_0 gnd vdd FILL
XFILL_4_1 gnd vdd FILL
XINVX1_17 opcode[1] gnd NOR2X1_2/B vdd INVX1
XNOR2X1_14 INVX4_1/A INVX2_7/Y gnd NOR2X1_14/Y vdd NOR2X1
XNOR2X1_36 NOR2X1_36/A INVX2_16/Y gnd INVX2_19/A vdd NOR2X1
XNAND3X1_14 NOR2X1_30/Y INVX4_1/Y INVX2_14/Y gnd NOR2X1_31/B vdd NAND3X1
XNOR2X1_25 A[1] B[1] gnd NOR2X1_41/A vdd NOR2X1
XOAI21X1_34 INVX2_10/Y INVX1_3/Y AOI21X1_14/Y gnd NOR2X1_13/B vdd OAI21X1
XFILL_4_0_1 gnd vdd FILL
XOAI21X1_23 B[5] A[5] INVX2_17/A gnd OAI21X1_24/C vdd OAI21X1
XOAI21X1_12 NAND2X1_9/Y NOR3X1_3/B INVX1_1/Y gnd INVX2_3/A vdd OAI21X1
XOAI21X1_45 XOR2X1_3/Y OR2X2_2/Y INVX1_15/Y gnd NOR2X1_28/A vdd OAI21X1
XFILL_4_2 gnd vdd FILL
XNOR2X1_15 OAI22X1_2/Y NOR2X1_15/B gnd NOR2X1_15/Y vdd NOR2X1
XNOR2X1_37 NOR2X1_33/A NOR2X1_42/A gnd INVX1_3/A vdd NOR2X1
XNAND3X1_15 NAND2X1_25/Y NAND2X1_26/Y OAI21X1_49/Y gnd NOR3X1_8/A vdd NAND3X1
XNOR2X1_26 B[2] A[2] gnd NOR2X1_26/Y vdd NOR2X1
XINVX1_18 opcode[0] gnd INVX1_18/Y vdd INVX1
XOAI21X1_35 NOR2X1_11/B INVX1_10/A INVX4_1/Y gnd NAND3X1_7/C vdd OAI21X1
XOAI21X1_46 INVX2_1/A NOR2X1_35/Y OAI21X1_2/B gnd AOI22X1_11/C vdd OAI21X1
XOAI21X1_24 INVX2_19/Y NAND2X1_14/Y OAI21X1_24/C gnd NOR3X1_2/A vdd OAI21X1
XOAI21X1_13 INVX2_3/A INVX2_2/A INVX2_7/A gnd OAI21X1_13/Y vdd OAI21X1
XFILL_4_3 gnd vdd FILL
XINVX1_19 opcode[3] gnd INVX1_19/Y vdd INVX1
XNOR2X1_38 NOR2X1_38/A NOR2X1_42/A gnd NOR2X1_38/Y vdd NOR2X1
XNAND3X1_16 NAND3X1_16/A NAND2X1_27/Y NAND3X1_16/C gnd NOR3X1_8/B vdd NAND3X1
XNOR2X1_16 INVX4_1/Y INVX2_7/Y gnd NAND3X1_8/B vdd NOR2X1
XFILL_2_1_0 gnd vdd FILL
XNOR2X1_27 B[3] A[3] gnd OAI22X1_4/D vdd NOR2X1
XFILL_7_0_0 gnd vdd FILL
XOAI21X1_47 OAI21X1_2/B INVX2_19/Y AOI22X1_12/Y gnd NOR2X1_39/A vdd OAI21X1
XOAI21X1_36 NOR2X1_9/B INVX2_9/A INVX2_14/Y gnd NAND3X1_6/C vdd OAI21X1
XOAI21X1_25 OAI21X1_25/A AOI21X1_8/Y NOR3X1_2/Y gnd OAI21X1_25/Y vdd OAI21X1
XOAI21X1_14 INVX1_2/Y INVX1_3/Y AOI22X1_6/Y gnd NOR2X1_7/B vdd OAI21X1
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XAND2X2_1 INVX1_19/Y opcode[2] gnd AND2X2_1/Y vdd AND2X2
XNOR2X1_17 opcode[0] opcode[1] gnd INVX2_18/A vdd NOR2X1
XNOR2X1_39 NOR2X1_39/A NOR2X1_39/B gnd NOR2X1_39/Y vdd NOR2X1
XNAND3X1_17 AOI22X1_2/D AND2X2_6/Y OR2X2_4/Y gnd NAND3X1_17/Y vdd NAND3X1
XNOR2X1_28 NOR2X1_28/A NOR2X1_28/B gnd NOR2X1_31/A vdd NOR2X1
XFILL_2_1_1 gnd vdd FILL
XFILL_2_1 gnd vdd FILL
XFILL_7_0_1 gnd vdd FILL
XOAI21X1_48 NOR2X1_31/Y OAI21X1_48/B NOR2X1_39/Y gnd BUFX2_3/A vdd OAI21X1
XOAI21X1_26 NOR2X1_31/A AOI21X1_7/C INVX2_9/Y gnd OAI21X1_26/Y vdd OAI21X1
XOAI21X1_37 AOI21X1_15/Y INVX1_7/A INVX2_14/A gnd NAND3X1_8/C vdd OAI21X1
XOAI21X1_15 INVX2_2/Y INVX2_5/Y AOI22X1_7/Y gnd NOR2X1_7/A vdd OAI21X1
XAND2X2_2 INVX2_6/A AND2X2_2/B gnd AND2X2_2/Y vdd AND2X2
XINVX1_2 A[5] gnd INVX1_2/Y vdd INVX1
XNOR2X1_18 INVX1_12/Y INVX2_10/Y gnd NOR2X1_20/B vdd NOR2X1
XNOR2X1_29 NOR2X1_23/Y INVX1_9/A gnd INVX2_14/A vdd NOR2X1
XNAND3X1_18 OAI21X1_50/Y NAND3X1_17/Y INVX2_7/A gnd NAND3X1_18/Y vdd NAND3X1
XFILL_2_2 gnd vdd FILL
XOAI21X1_38 INVX1_13/Y INVX2_11/Y NAND3X1_8/C gnd OAI21X1_38/Y vdd OAI21X1
XOAI21X1_49 A[1] B[1] INVX2_17/A gnd OAI21X1_49/Y vdd OAI21X1
XOAI21X1_27 NOR2X1_28/B NOR2X1_28/A NOR2X1_30/Y gnd OAI21X1_27/Y vdd OAI21X1
XOAI21X1_16 NOR2X1_6/Y OAI21X1_13/Y NOR2X1_7/Y gnd NOR2X1_8/B vdd OAI21X1
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XOR2X2_1 B[3] A[3] gnd OR2X2_1/Y vdd OR2X2
XNOR2X1_19 B[7] A[7] gnd NOR2X1_20/A vdd NOR2X1
XFILL_5_1_0 gnd vdd FILL
XAND2X2_3 A[1] B[1] gnd AND2X2_3/Y vdd AND2X2
XFILL_2_3 gnd vdd FILL
XOAI22X1_1 INVX2_19/Y INVX1_9/Y NOR2X1_23/Y INVX2_17/Y gnd NOR2X1_13/A vdd OAI22X1
XNAND2X1_30 B[0] INVX2_15/Y gnd NOR2X1_43/A vdd NAND2X1
XINVX2_10 A[7] gnd INVX2_10/Y vdd INVX2
XOAI21X1_39 INVX2_11/Y NAND2X1_2/Y AOI22X1_10/Y gnd NOR2X1_15/B vdd OAI21X1
XOAI21X1_17 NOR2X1_31/A INVX2_2/A AND2X2_2/Y gnd AOI21X1_10/A vdd OAI21X1
XOAI21X1_28 INVX2_14/Y OAI21X1_26/Y NOR2X1_11/Y gnd NAND3X1_5/A vdd OAI21X1
XFILL_5_1_1 gnd vdd FILL
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XOR2X2_2 OR2X2_2/A B[2] gnd OR2X2_2/Y vdd OR2X2
XNAND2X1_20 opcode[0] opcode[1] gnd NOR2X1_33/A vdd NAND2X1
XNAND2X1_31 A[1] B[1] gnd AOI22X1_2/D vdd NAND2X1
XAND2X2_4 B[2] A[2] gnd NOR2X1_5/A vdd AND2X2
XOAI22X1_2 INVX2_17/Y NOR2X1_20/A INVX4_1/Y INVX2_5/Y gnd OAI22X1_2/Y vdd OAI22X1
XINVX2_11 A[6] gnd INVX2_11/Y vdd INVX2
XOAI21X1_29 INVX2_6/Y INVX1_4/A NAND2X1_14/Y gnd INVX1_7/A vdd OAI21X1
XOAI21X1_18 AOI22X1_2/Y NOR2X1_3/Y AOI22X1_8/Y gnd AOI21X1_7/B vdd OAI21X1
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XOR2X2_3 OR2X2_3/A B[1] gnd OR2X2_3/Y vdd OR2X2
.ends

